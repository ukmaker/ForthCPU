library verilog;
use verilog.vl_types.all;
entity ts_dgflow_fsm is
    generic(
        st_idle_d       : integer := 0;
        st_load_offsets_d: integer := 1;
        st_toffset_1_d  : integer := 3;
        st_read_vbe1_d  : integer := 2;
        st_wait_vbe2_d  : integer := 6;
        st_read_vbe2_d  : integer := 4;
        st_wait_vbe3_d  : integer := 5;
        st_read_vbe3_d  : integer := 7;
        st_delvbe1_d    : integer := 15;
        st_delvbe2_d    : integer := 14;
        st_mul_x_2_d    : integer := 12;
        st_y_from_2x_add_x_d: integer := 13;
        st_mul_y_d      : integer := 9;
        st_wait_mul_y_d : integer := 11;
        st_mul_y_done_d : integer := 10;
        st_mul_x_d      : integer := 8;
        st_wait_mul_x_d : integer := 24;
        st_mul_x_done_d : integer := 28;
        st_diff_ydelta_xdelta_d: integer := 30;
        st_rshift_15_d  : integer := 31;
        st_tout_kelvin_d: integer := 29;
        st_tout_dec_d   : integer := 25;
        st_read_pre_ave_d: integer := 17;
        st_mul_const_d  : integer := 19;
        st_wait_mul_const_d: integer := 18;
        st_mul_const_done_d: integer := 22;
        st_add_tmeas_ave_d: integer := 23;
        st_lshift_3_d   : integer := 21;
        st_lshift_4_d   : integer := 20;
        st_store_tmeas_d: integer := 16;
        st_done_d       : integer := 26
    );
    port(
        asc_clk         : in     vl_logic;
        ts_resetb       : in     vl_logic;
        ts_start_dgflow : in     vl_logic;
        ts_cic_data_ready: in     vl_logic;
        ts_ave_en       : in     vl_logic;
        ts_ave_8        : in     vl_logic;
        ts_first_ave_flag: in     vl_logic;
        ts_pre_ave_zero : in     vl_logic;
        ts_mon_data_valid: out    vl_logic;
        ts_start_mul    : out    vl_logic;
        ts_clr_acc_reg  : out    vl_logic;
        ts_rshift_acc_reg_from_dgflow: out    vl_logic;
        ts_mul_done     : in     vl_logic;
        ts_ld_from_alu_tmeas_reg: out    vl_logic;
        ts_ld_from_alu_toffset_reg: out    vl_logic;
        ts_ld_from_alu_vbe_diff_reg: out    vl_logic;
        ts_ld_from_alu_prod_vbe_diff_reg: out    vl_logic;
        ts_rd_from_alu_m_filter_reg: out    vl_logic;
        ts_rd_from_alu_m_x_reg: out    vl_logic;
        ts_rd_from_alu_m_273: out    vl_logic;
        ts_rd_from_alu_m_trim_reg: out    vl_logic;
        ts_rd_from_alu_m_tmeas_reg: out    vl_logic;
        ts_rd_from_alu_m_toffset_reg: out    vl_logic;
        ts_rd_from_alu_m_vbe_diff_reg: out    vl_logic;
        ts_rd_from_alu_m_prod_datain: out    vl_logic;
        ts_rd_from_alu_m_acc: out    vl_logic;
        ts_rd_from_alu_acc_vbe_diff_reg: out    vl_logic;
        ts_rd_from_alu_acc_selfheat_reg: out    vl_logic;
        ts_rd_from_alu_acc_filter_reg: out    vl_logic;
        ts_rd_from_alu_acc_datain: out    vl_logic;
        ts_rd_from_alu_acc_prod_datain: out    vl_logic;
        ts_rd_from_alu_acc_x_reg: out    vl_logic;
        ts_rd_from_alu_acc_m: out    vl_logic;
        ts_rd_from_alu_acc_q: out    vl_logic;
        ts_rd_from_alu_q_filter_reg: out    vl_logic;
        ts_rd_from_alu_q_vbe_diff_reg: out    vl_logic;
        ts_rd_from_alu_q_datain: out    vl_logic;
        ts_rd_from_alu_q_ave_reg: out    vl_logic;
        alu_mode        : out    vl_logic_vector(2 downto 0);
        ts_dgflow_done_clr: in     vl_logic;
        ts_dgflow_done  : out    vl_logic;
        ts_dgflow_done_reg: out    vl_logic;
        ts_disable_cal_tst: in     vl_logic
    );
end ts_dgflow_fsm;
