library verilog;
use verilog.vl_types.all;
entity cfg_pdrv is
    generic(
        FLASH_MEM       : integer := 1
    );
    port(
        spi2nd_men      : out    vl_logic;
        p16_in          : out    vl_logic_vector(15 downto 0);
        extspi_out      : out    vl_logic;
        persist_out_cib : out    vl_logic_vector(15 downto 0);
        data_o_1st      : out    vl_logic_vector(15 downto 0);
        data_oe_1st     : out    vl_logic_vector(15 downto 0);
        mcsn_o_1st      : out    vl_logic_vector(7 downto 0);
        mcsn_oe_1st     : out    vl_logic_vector(7 downto 0);
        mclk_o_1st      : out    vl_logic;
        mclk_oe_1st     : out    vl_logic;
        mclk_byp_o      : out    vl_logic;
        mclk_byp_oe     : out    vl_logic;
        docson_o        : out    vl_logic;
        docson_oe       : out    vl_logic;
        busy_o_1st      : out    vl_logic;
        busy_oe_1st     : out    vl_logic;
        initn_o         : out    vl_logic;
        initn_oe        : out    vl_logic;
        donep_o         : out    vl_logic;
        donep_oe        : out    vl_logic;
        int_spi_mclk    : out    vl_logic;
        int_spi_data    : out    vl_logic_vector(15 downto 0);
        int_spi_mcsn    : out    vl_logic_vector(7 downto 0);
        cfgmode_cfg     : out    vl_logic;
        spi2nd_miso_i   : out    vl_logic;
        INT_SPI_CTRL    : in     vl_logic_vector(1 downto 0);
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        programn_tog    : in     vl_logic;
        tck_pin         : in     vl_logic;
        tdi             : in     vl_logic;
        cclk_in         : in     vl_logic;
        sspi_si         : in     vl_logic;
        din_16          : in     vl_logic_vector(15 downto 0);
        miso_i_2nd      : in     vl_logic;
        ctrl_cpol       : in     vl_logic;
        ctrl_done_opt   : in     vl_logic_vector(1 downto 0);
        ctrl_initn_opt  : in     vl_logic_vector(1 downto 0);
        ref_boot0       : in     vl_logic;
        ref_boot1       : in     vl_logic;
        ref_boot2       : in     vl_logic;
        initn_tmr       : in     vl_logic;
        goe_tmr         : in     vl_logic;
        done_tmr        : in     vl_logic;
        isc_operational : in     vl_logic;
        njbse_bypass    : in     vl_logic;
        njbse_fthrough  : in     vl_logic;
        cfg_mclk_o      : in     vl_logic;
        cfg_mclk_oe     : in     vl_logic;
        cfg_mclk_byp_o  : in     vl_logic;
        cfg_mclk_byp_oe : in     vl_logic;
        cfg_data_o      : in     vl_logic_vector(15 downto 0);
        cfg_data_oe     : in     vl_logic_vector(15 downto 0);
        cfg_mcsn_o      : in     vl_logic_vector(7 downto 0);
        cfg_mcsn_oe     : in     vl_logic_vector(7 downto 0);
        cfg_sd_out      : in     vl_logic;
        cfg_busy_o      : in     vl_logic;
        cfg_busy_oe     : in     vl_logic;
        shiftdr_ss      : in     vl_logic;
        ShiftDR         : in     vl_logic;
        jpspi_en_norm   : in     vl_logic;
        jpspi_en_stack  : in     vl_logic;
        jpspi_en_int    : in     vl_logic;
        jpspi_param     : in     vl_logic_vector(7 downto 0);
        njshf_dat0      : in     vl_logic;
        njshf_dat_nd    : in     vl_logic;
        njpspi_en_norm  : in     vl_logic;
        njpspi_en_stack : in     vl_logic;
        njpspi_en_int   : in     vl_logic;
        njpspi_param    : in     vl_logic_vector(7 downto 0);
        spi2nd_cfg_mcsn : in     vl_logic;
        spi2nd_cfg_mcsn_2d: in     vl_logic;
        spi2nd_mclk_o   : in     vl_logic;
        spi2nd_mclk_oe  : in     vl_logic;
        spi2nd_mosi_o   : in     vl_logic;
        spi2nd_mosi_oe  : in     vl_logic;
        int_spi_din     : in     vl_logic_vector(15 downto 0);
        mc1_persist_cap : in     vl_logic;
        fsd_persist_initn: in     vl_logic;
        fsd_persist_done: in     vl_logic;
        cib_persist_in  : in     vl_logic_vector(15 downto 0);
        persist_slave   : in     vl_logic
    );
end cfg_pdrv;
