library verilog;
use verilog.vl_types.all;
entity jtag_cntl is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 1;
        DECRYPTION      : integer := 1
    );
    port(
        tlreset         : out    vl_logic;
        rti             : out    vl_logic;
        ShiftDR         : out    vl_logic;
        UpdateDR        : out    vl_logic;
        CaptureDR       : out    vl_logic;
        ClockIR         : out    vl_logic;
        ClockDR         : out    vl_logic;
        ShiftIR         : out    vl_logic;
        UpdateIR        : out    vl_logic;
        CaptureIR       : out    vl_logic;
        upir_ss         : out    vl_logic;
        selir_ss        : out    vl_logic;
        updr_ss         : out    vl_logic;
        seldr_ss        : out    vl_logic;
        shiftdr_ss      : out    vl_logic;
        capdr_ss_r      : out    vl_logic;
        rti_r           : out    vl_logic;
        upir_ss_r       : out    vl_logic;
        exit1dr_ss_r    : out    vl_logic;
        isc_data_shift_iq: out    vl_logic;
        isc_addr_shift_iq: out    vl_logic;
        verify_id_iq    : out    vl_logic;
        idcode_pub_iq   : out    vl_logic;
        uidcode_pub_iq  : out    vl_logic;
        usercode_iq     : out    vl_logic;
        read_temp_iq    : out    vl_logic;
        lsc_device_ctrl_iq: out    vl_logic;
        lsc_shift_password_iq: out    vl_logic;
        lsc_read_status_mq: out    vl_logic;
        lsc_read_mfg_status_mq: out    vl_logic;
        lsc_refresh_iq  : out    vl_logic;
        lsc_bitstream_burst_iq: out    vl_logic;
        idcode_prv_iq   : out    vl_logic;
        lsc_read_pes_mq : out    vl_logic;
        lsc_prog_ctrl0_iq: out    vl_logic;
        lsc_read_ctrl0_iq: out    vl_logic;
        lsc_reset_crc_iq: out    vl_logic;
        lsc_read_crc_iq : out    vl_logic;
        lsc_write_comp_dic_iq: out    vl_logic;
        lsc_read_comp_dic_mq: out    vl_logic;
        sf_prog_ucode_iq: out    vl_logic;
        sf_program_iq   : out    vl_logic;
        sf_read_iq      : out    vl_logic;
        sf_erase_iq     : out    vl_logic;
        sf_prog_done_iq : out    vl_logic;
        sf_erase_done_iq: out    vl_logic;
        sf_prog_sec_iq  : out    vl_logic;
        sf_init_addr_iq : out    vl_logic;
        sf_write_addr_iq: out    vl_logic;
        sf_prog_incr_rti_iq: out    vl_logic;
        sf_prog_incr_enc_iq: out    vl_logic;
        sf_prog_incr_cmp_iq: out    vl_logic;
        sf_prog_incr_cne_iq: out    vl_logic;
        sf_vfy_incr_rti_iq: out    vl_logic;
        sf_prog_sed_crc_iq: out    vl_logic;
        sf_read_sed_crc_iq: out    vl_logic;
        sf_write_bus_addr_iq: out    vl_logic;
        sf_pcs_write_iq : out    vl_logic;
        sf_pcs_read_iq  : out    vl_logic;
        sf_ebr_write_iq : out    vl_logic;
        sf_ebr_read_iq  : out    vl_logic;
        fl_prog_ucode_iq: out    vl_logic;
        fl_erase_iq     : out    vl_logic;
        fl_prog_done_iq : out    vl_logic;
        fl_prog_sec_iq  : out    vl_logic;
        fl_prog_secplus_iq: out    vl_logic;
        fl_init_addr_iq : out    vl_logic;
        fl_write_addr_iq: out    vl_logic;
        fl_prog_incr_nv_iq: out    vl_logic;
        fl_read_incr_nv_iq: out    vl_logic;
        fl_prog_password_iq: out    vl_logic;
        fl_read_password_iq: out    vl_logic;
        fl_prog_cipher_key_iq: out    vl_logic;
        fl_read_cipher_key_iq: out    vl_logic;
        fl_prog_feature_iq: out    vl_logic;
        fl_read_feature_iq: out    vl_logic;
        fl_prog_feabits_iq: out    vl_logic;
        fl_read_feabits_iq: out    vl_logic;
        fl_prog_otps_iq : out    vl_logic;
        fl_read_otps_iq : out    vl_logic;
        fl_init_addr_ufm_iq: out    vl_logic;
        fl_erase_tag_iq : out    vl_logic;
        fl_prog_tag_iq  : out    vl_logic;
        fl_read_tag_iq  : out    vl_logic;
        fl_prog_pes_mq  : out    vl_logic;
        fl_prog_trim_mq : out    vl_logic;
        fl_prog_mes_mq  : out    vl_logic;
        fl_prog_hes_mq  : out    vl_logic;
        fl_read_trim_mq : out    vl_logic;
        fl_read_mes_mq  : out    vl_logic;
        fl_read_hes_mq  : out    vl_logic;
        ef_init_addr_iq : out    vl_logic;
        ef_write_addr_iq: out    vl_logic;
        ef_prog_password_iq: out    vl_logic;
        ef_read_password_iq: out    vl_logic;
        ef_prog_cipher_key_iq: out    vl_logic;
        ef_read_cipher_key_iq: out    vl_logic;
        ef_prog_feature_iq: out    vl_logic;
        ef_read_feature_iq: out    vl_logic;
        ef_prog_feabits_iq: out    vl_logic;
        ef_read_feabits_iq: out    vl_logic;
        ef_prog_otps_iq : out    vl_logic;
        ef_read_otps_iq : out    vl_logic;
        ef_prog_pes_mq  : out    vl_logic;
        ef_prog_trim_mq : out    vl_logic;
        ef_prog_mes_mq  : out    vl_logic;
        ef_prog_hes_mq  : out    vl_logic;
        ef_read_trim_mq : out    vl_logic;
        ef_read_mes_mq  : out    vl_logic;
        ef_read_hes_mq  : out    vl_logic;
        ef_prog_main_rmr_mq: out    vl_logic;
        ef_prog_efrtest_mq: out    vl_logic;
        ef_prog_efctest_mq: out    vl_logic;
        ef_prog_efarray_mq: out    vl_logic;
        ef_read_efrtest_mq: out    vl_logic;
        ef_read_efctest_mq: out    vl_logic;
        ef_read_efarray_mq: out    vl_logic;
        mfg_mtest_mq    : out    vl_logic;
        mfg_mtrim_mq    : out    vl_logic;
        mfg_mdata_mq    : out    vl_logic;
        lsc_i2ci_crbr_wt_iq: out    vl_logic;
        lsc_i2ci_txdr_wt_iq: out    vl_logic;
        lsc_i2ci_rxdr_rd_iq: out    vl_logic;
        lsc_i2ci_sr_rd_iq: out    vl_logic;
        isptcy_ener1    : out    vl_logic;
        isptcy_ener2    : out    vl_logic;
        isptcy_resetb   : out    vl_logic;
        isptcy_shcap    : out    vl_logic;
        isptcy_update   : out    vl_logic;
        isptcy_rtier1   : out    vl_logic;
        isptcy_rtier2   : out    vl_logic;
        isptcy_tdi      : out    vl_logic;
        bsrclk          : out    vl_logic;
        shiftdr_bs      : out    vl_logic;
        updatedr_bs     : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        bsmode_pcs      : out    vl_logic;
        ac_mode         : out    vl_logic;
        ac_clear        : out    vl_logic;
        ac_test         : out    vl_logic;
        tsall_ctrl      : out    vl_logic;
        isc_test_mode   : out    vl_logic;
        isc_enabled     : out    vl_logic;
        isc_disable_completing: out    vl_logic;
        jaccess_sram    : out    vl_logic;
        jaccess_flash   : out    vl_logic;
        jaccess_fl_norm : out    vl_logic;
        jaccess_fl_sudo : out    vl_logic;
        jaccess_fl_safe : out    vl_logic;
        jaccess_efuse   : out    vl_logic;
        jaccess_ef_norm : out    vl_logic;
        jaccess_ef_sudo : out    vl_logic;
        jaccess_ef_safe : out    vl_logic;
        jaccess_tag     : out    vl_logic;
        jaccess_flash_all: out    vl_logic;
        jenable_offl    : out    vl_logic;
        mfg_dat         : out    vl_logic_vector(119 downto 0);
        mfg_en          : out    vl_logic;
        rti2d           : out    vl_logic;
        jconfig_dat     : out    vl_logic_vector(3 downto 0);
        jsector_dat     : out    vl_logic_vector(7 downto 0);
        jbuf128_dat     : out    vl_logic_vector(127 downto 0);
        jbuf8_dat       : out    vl_logic_vector(7 downto 0);
        jbuf8_rdy       : out    vl_logic;
        tdrclk_sw_i     : out    vl_logic;
        jexit_fl_offline: out    vl_logic;
        jexit_normal    : out    vl_logic;
        j_enable_qual   : out    vl_logic;
        j_enable_x_qual : out    vl_logic;
        j_disable_qual  : out    vl_logic;
        jrst_isc_done_i : out    vl_logic;
        jset_isc_done_i : out    vl_logic;
        jtag_active     : out    vl_logic;
        jsec_dsr        : out    vl_logic;
        tdo_out         : out    vl_logic;
        tdo_oe_out      : out    vl_logic;
        tdi_sram_asr    : out    vl_logic;
        tdi_bscan       : out    vl_logic;
        tdi_rmr         : out    vl_logic;
        tdi_iscan       : out    vl_logic;
        jsel_bsr        : out    vl_logic;
        jsel_sram_asr   : out    vl_logic;
        jsel_rmr        : out    vl_logic;
        ins_dsr_1bit    : out    vl_logic;
        ins_dsr_1byte   : out    vl_logic;
        tdi_dsr_1bit    : out    vl_logic;
        tdi_dsr_1byte   : out    vl_logic_vector(7 downto 0);
        jburst_pause    : out    vl_logic;
        jburst_01       : out    vl_logic;
        jburst_08       : out    vl_logic;
        j_ins_prog_com  : out    vl_logic;
        jburst_en       : out    vl_logic;
        jpspi_en_norm   : out    vl_logic;
        jpspi_en_stack  : out    vl_logic;
        jpspi_en_int    : out    vl_logic;
        jpspi_param     : out    vl_logic_vector(7 downto 0);
        iscan_en        : out    vl_logic_vector(7 downto 0);
        mfg_scan_test_mode: out    vl_logic;
        por             : in     vl_logic;
        tck             : in     vl_logic;
        tdi             : in     vl_logic;
        tms             : in     vl_logic;
        busy_seldr      : in     vl_logic;
        isc_done        : in     vl_logic;
        j_com_word4_dat : in     vl_logic_vector(127 downto 0);
        jinstr_cap      : in     vl_logic_vector(7 downto 0);
        jconfig_cap     : in     vl_logic_vector(7 downto 0);
        ctrl_tran_edit  : in     vl_logic;
        mfg_prog_sel    : in     vl_logic_vector(3 downto 0);
        mfg_iscan_sel   : in     vl_logic_vector(2 downto 0);
        mfg_iscan_en    : in     vl_logic;
        mfg_pshf_sel    : in     vl_logic;
        mfg_tckrti      : in     vl_logic;
        dsr_out_jtag    : in     vl_logic;
        sram_asr_out    : in     vl_logic;
        p8_in           : in     vl_logic_vector(7 downto 0);
        bscan_out       : in     vl_logic;
        isptracy_er1_out: in     vl_logic;
        isptracy_er2_out: in     vl_logic;
        rmr_dout        : in     vl_logic;
        iscan_out       : in     vl_logic_vector(7 downto 0);
        extspi_out      : in     vl_logic;
        mc1_er1_exist   : in     vl_logic;
        mc1_er2_exist   : in     vl_logic;
        scan_test_mode  : in     vl_logic;
        mc1_scan_test_en: in     vl_logic_vector(3 downto 0);
        stm_tap_state   : in     vl_logic_vector(3 downto 0)
    );
end jtag_cntl;
