library verilog;
use verilog.vl_types.all;
entity reno_dig_io is
    generic(
        MCLK_8MHZ_PERIOD: integer := 125
    );
    port(
        fsafeb          : out    vl_logic;
        ana_rst_b       : in     vl_logic;
        wrclk_in        : in     vl_logic;
        clk_loss_off    : in     vl_logic;
        wrclk_lost      : out    vl_logic;
        por_off         : in     vl_logic;
        por_n           : out    vl_logic;
        resetb          : inout  vl_logic;
        resetb_in_pin   : out    vl_logic;
        resetb_out_pin  : in     vl_logic;
        mclkout         : out    vl_logic;
        rst_osc_b       : in     vl_logic;
        rst_osc_tmr_b   : in     vl_logic;
        mclk            : in     vl_logic;
        rst_abg_b       : in     vl_logic;
        bg_caldone      : out    vl_logic;
        dac_resetb      : in     vl_logic;
        dac_ready       : out    vl_logic;
        sda             : inout  vl_logic;
        scl             : in     vl_logic;
        sda_out         : in     vl_logic;
        sda_in          : out    vl_logic;
        scl_in          : out    vl_logic;
        i2cdet_compout  : out    vl_logic;
        i2cdet_clk      : in     vl_logic;
        i2cdet_resetb   : in     vl_logic;
        i2cdet_tapsel   : in     vl_logic_vector(2 downto 0);
        gpio_1          : inout  vl_logic;
        gpio_2          : inout  vl_logic;
        gpio_3          : inout  vl_logic;
        gpio_4          : inout  vl_logic;
        gpio_5          : inout  vl_logic;
        gpio_6          : inout  vl_logic;
        gpio_7          : inout  vl_logic;
        gpio_8          : inout  vl_logic;
        gpio_9          : inout  vl_logic;
        gpio_10         : inout  vl_logic;
        wgpio_1         : in     vl_logic;
        wgpio_2         : in     vl_logic;
        wgpio_3         : in     vl_logic;
        wgpio_4         : in     vl_logic;
        wgpio_5         : in     vl_logic;
        wgpio_6         : in     vl_logic;
        wgpio_7         : in     vl_logic;
        wgpio_8         : in     vl_logic;
        wgpio_9         : in     vl_logic;
        wgpio_10        : in     vl_logic;
        rgpio_1         : out    vl_logic;
        rgpio_2         : out    vl_logic;
        rgpio_3         : out    vl_logic;
        rgpio_4         : out    vl_logic;
        rgpio_5         : out    vl_logic;
        rgpio_6         : out    vl_logic;
        rgpio_7         : out    vl_logic;
        rgpio_8         : out    vl_logic;
        rgpio_9         : out    vl_logic;
        rgpio_10        : out    vl_logic;
        gpio_oeb        : in     vl_logic_vector(9 downto 0);
        gpio_pldn_en    : in     vl_logic_vector(9 downto 0);
        cfg_vm          : inout  vl_logic_vector(7 downto 0);
        ldshdwreg       : in     vl_logic;
        ldmshdw         : in     vl_logic;
        ldsshdw         : in     vl_logic;
        rdshdw          : in     vl_logic;
        reset_in_b      : in     vl_logic
    );
end reno_dig_io;
