library verilog;
use verilog.vl_types.all;
entity config_plus is
    port(
        int_csspi0n     : out    vl_logic;
        int_mclk        : out    vl_logic;
        int_sispi       : out    vl_logic;
        sci_initen      : out    vl_logic_vector(1 downto 0);
        sci_rst_n       : out    vl_logic;
        ss_addr         : out    vl_logic_vector(7 downto 0);
        ss_clk          : out    vl_logic;
        ss_rst          : out    vl_logic;
        ss_stb          : out    vl_logic;
        ss_wdata        : out    vl_logic_vector(7 downto 0);
        ss_we           : out    vl_logic;
        bsrclk          : out    vl_logic;
        bsrtdi          : out    vl_logic;
        bsmode          : out    vl_logic;
        intest          : out    vl_logic;
        shbsrn          : out    vl_logic;
        treset          : out    vl_logic;
        ts_all          : out    vl_logic;
        updtbsr         : out    vl_logic;
        addr_clk        : out    vl_logic;
        asr_addr_in     : out    vl_logic;
        asr_en_addr     : out    vl_logic;
        asr_en_incr     : out    vl_logic;
        asr_init_0      : out    vl_logic;
        asr_shift_1st   : out    vl_logic;
        asr_shift_2nd   : out    vl_logic;
        asr_shift_3rd   : out    vl_logic;
        bg_trim         : out    vl_logic_vector(15 downto 0);
        bgoff           : out    vl_logic;
        cfg_addr_slew   : out    vl_logic;
        cfg_addr_por_n  : out    vl_logic;
        cfg_data_cap    : out    vl_logic;
        cfg_data_flt    : out    vl_logic;
        cfg_data_por_n  : out    vl_logic;
        cfg_data_pre    : out    vl_logic;
        cfg_data_wr     : out    vl_logic;
        data_clk        : out    vl_logic;
        dsr_cfg_d       : out    vl_logic_vector(63 downto 0);
        dsr_got_data    : out    vl_logic;
        dsr_ld_rdbkd    : out    vl_logic;
        dsr_reset_n     : out    vl_logic;
        dsr_shift_d     : out    vl_logic_vector(1 downto 0);
        dtr_clk         : out    vl_logic;
        dtr_instr       : out    vl_logic;
        dtr_start       : out    vl_logic;
        mfg_bits        : out    vl_logic_vector(47 downto 0);
        osc_dis         : out    vl_logic;
        osc_ena         : out    vl_logic;
        osc_trim        : out    vl_logic_vector(7 downto 0);
        poroff          : out    vl_logic;
        sram_ppt_addr   : out    vl_logic_vector(3 downto 0);
        trim_bits       : out    vl_logic_vector(63 downto 0);
        csspin          : out    vl_logic;
        init_n          : out    vl_logic;
        mclk_out        : out    vl_logic;
        pad_done        : out    vl_logic;
        scl             : out    vl_logic;
        sda             : out    vl_logic;
        si              : out    vl_logic;
        so              : out    vl_logic;
        tdo             : out    vl_logic;
        done_md_n       : out    vl_logic;
        done_ts         : out    vl_logic;
        init_md_n       : out    vl_logic;
        init_ts         : out    vl_logic;
        i2c_md_n        : out    vl_logic;
        jtag_md_n       : out    vl_logic;
        mclk_ts         : out    vl_logic;
        mspi_md_n       : out    vl_logic;
        pll_mfg_ts      : out    vl_logic_vector(1 downto 0);
        pll_mfg_md_n    : out    vl_logic_vector(1 downto 0);
        program_md_n    : out    vl_logic;
        scl_ts          : out    vl_logic;
        sda_ts          : out    vl_logic;
        si_md_n         : out    vl_logic;
        si_ts           : out    vl_logic;
        so_md_n         : out    vl_logic;
        so_ts           : out    vl_logic;
        tdo_ts          : out    vl_logic;
        done_goe        : out    vl_logic;
        done_gwe        : out    vl_logic;
        freeze_io       : out    vl_logic;
        freeze_mib      : out    vl_logic;
        gsrn            : out    vl_logic;
        por_n           : out    vl_logic;
        cib_i2c_scl     : out    vl_logic;
        cib_i2c_sclen   : out    vl_logic;
        cib_i2c_sda     : out    vl_logic;
        cib_i2c_sdaen   : out    vl_logic;
        cib_mspi_csn    : out    vl_logic_vector(7 downto 1);
        jce             : out    vl_logic_vector(2 downto 1);
        jrstn           : out    vl_logic;
        jrti            : out    vl_logic_vector(2 downto 1);
        jshift          : out    vl_logic;
        jtck            : out    vl_logic;
        jtdi            : out    vl_logic;
        jupdate         : out    vl_logic;
        auto_done       : out    vl_logic;
        cib_done        : out    vl_logic;
        cib_freeze_io   : out    vl_logic;
        cib_last_addr   : out    vl_logic_vector(7 downto 0);
        sflag           : out    vl_logic;
        stdby           : out    vl_logic;
        stop            : out    vl_logic;
        usrclk_cib      : out    vl_logic;
        sed_clk_out     : out    vl_logic;
        sed_done        : out    vl_logic;
        sed_inprog      : out    vl_logic;
        sed_err         : out    vl_logic;
        es_o            : out    vl_logic_vector(35 downto 0);
        fl_row          : out    vl_logic_vector(14 downto 0);
        fl_ufm_row_sel_all: out    vl_logic;
        fl_ufm_row_sel_none: out    vl_logic;
        fl_cfg_row_sel_all: out    vl_logic;
        fl_cfg_row_sel_none: out    vl_logic;
        fl_trim_row_sel_all: out    vl_logic;
        fl_trim_row_sel_none: out    vl_logic;
        fl_feat_row_sel_all: out    vl_logic;
        fl_feat_row_sel_none: out    vl_logic;
        fl_era_ufm      : out    vl_logic;
        fl_era_cfg      : out    vl_logic;
        fl_era_trim     : out    vl_logic;
        fl_era_feat     : out    vl_logic;
        fl_prg_ufm      : out    vl_logic;
        fl_prg_cfg      : out    vl_logic;
        fl_prg_tf       : out    vl_logic;
        fl_read_ufm     : out    vl_logic;
        fl_read_cfg     : out    vl_logic;
        fl_read_tf      : out    vl_logic;
        fl_erase_setup  : out    vl_logic;
        fl_erapdis      : out    vl_logic;
        fl_erase_pulse  : out    vl_logic;
        fl_pwtc_well    : out    vl_logic;
        fl_prg_pulse    : out    vl_logic_vector(3 downto 0);
        fl_prog_disch   : out    vl_logic;
        fl_prg_pwtc     : out    vl_logic;
        fl_en_vreg_mon  : out    vl_logic;
        fl_era_ver      : out    vl_logic;
        fl_scp          : out    vl_logic;
        fl_softprg      : out    vl_logic;
        fl_verify       : out    vl_logic;
        fl_flash_en     : out    vl_logic;
        fl_reg_enable   : out    vl_logic;
        fl_subrow_mvena_ufm: out    vl_logic;
        fl_subrow_mvenall_ufm: out    vl_logic;
        fl_subrow_hvena_ufm: out    vl_logic;
        fl_subrow_hvenall_ufm: out    vl_logic;
        fl_subrow_mvena_cfg: out    vl_logic;
        fl_subrow_mvenall_cfg: out    vl_logic;
        fl_subrow_hvena_cfg: out    vl_logic;
        fl_subrow_hvenall_cfg: out    vl_logic;
        fl_subrow_mvena_tf: out    vl_logic;
        fl_subrow_hvena_tf: out    vl_logic;
        fl_sa_enall     : out    vl_logic;
        fl_sa_ena       : out    vl_logic;
        fl_prgdrv_enall : out    vl_logic;
        fl_prgdrv_ena   : out    vl_logic;
        fl_col_shift    : out    vl_logic;
        fl_colstart     : out    vl_logic_vector(3 downto 0);
        fl_col_rst      : out    vl_logic;
        fl_readpart     : out    vl_logic_vector(3 downto 0);
        fl_wor_eval     : out    vl_logic;
        fl_wand_eval    : out    vl_logic;
        fl_capture_dout : out    vl_logic;
        fl_src_clamp    : out    vl_logic;
        fl_scpv         : out    vl_logic;
        fl_drain_ctrl   : out    vl_logic;
        fl_sel_6p5v     : out    vl_logic;
        fl_prestep_in_neg: out    vl_logic_vector(2 downto 0);
        fl_step_in_neg  : out    vl_logic_vector(2 downto 0);
        fl_ppt_en       : out    vl_logic;
        fl_ppt_pset     : out    vl_logic;
        fl_ppt_rowsel   : out    vl_logic;
        fl_ready_rst    : out    vl_logic;
        fl_mfg_margin_en: out    vl_logic;
        flash_clk_mfg   : out    vl_logic;
        mux32_out1_mfg  : out    vl_logic;
        mux32_out2_mfg  : out    vl_logic;
        cfg_se          : out    vl_logic;
        sel_scan2       : out    vl_logic;
        i2cgcdr_1st     : out    vl_logic_vector(7 downto 0);
        i2cgcdr_2nd     : out    vl_logic_vector(7 downto 0);
        i2crxdr_1st     : out    vl_logic_vector(7 downto 0);
        i2crxdr_2nd     : out    vl_logic_vector(7 downto 0);
        i2csr_1st       : out    vl_logic_vector(7 downto 0);
        i2csr_2nd       : out    vl_logic_vector(7 downto 0);
        spirxdr         : out    vl_logic_vector(7 downto 0);
        spisr           : out    vl_logic_vector(7 downto 0);
        wbcrxdr         : out    vl_logic_vector(7 downto 0);
        wbcsr           : out    vl_logic_vector(7 downto 0);
        asr_length      : in     vl_logic_vector(13 downto 0);
        chipid          : in     vl_logic_vector(7 downto 0);
        device          : in     vl_logic_vector(2 downto 0);
        dsr_length      : in     vl_logic_vector(15 downto 0);
        idcode          : in     vl_logic_vector(31 downto 0);
        int_spid0       : in     vl_logic;
        bsout           : in     vl_logic;
        ss_ack          : in     vl_logic;
        ss_rdata        : in     vl_logic_vector(7 downto 0);
        asr_addr_out    : in     vl_logic;
        bg_cmp_out      : in     vl_logic;
        bg_stable       : in     vl_logic;
        cfg_osc         : in     vl_logic;
        dtr_out         : in     vl_logic_vector(31 downto 0);
        dsr_rdbk_dout   : in     vl_logic_vector(7 downto 0);
        proc_ring_osc   : in     vl_logic;
        pwrup_pur_n     : in     vl_logic;
        cclkin          : in     vl_logic;
        donein          : in     vl_logic;
        initin_n        : in     vl_logic;
        jtagenb         : in     vl_logic;
        pi_mcsn         : in     vl_logic;
        pfsafe          : in     vl_logic;
        programn        : in     vl_logic;
        pi_scl          : in     vl_logic;
        pi_sda          : in     vl_logic;
        pi_si           : in     vl_logic;
        pi_sn           : in     vl_logic;
        pi_so           : in     vl_logic;
        tck             : in     vl_logic;
        tdi             : in     vl_logic;
        tms             : in     vl_logic;
        mc1_auto_sel    : in     vl_logic;
        mc1_bl_float    : in     vl_logic;
        mc1_bypass_timer: in     vl_logic;
        mc1_clk_sel     : in     vl_logic;
        mc1_dis_bg      : in     vl_logic_vector(1 downto 0);
        mc1_dis_osc     : in     vl_logic;
        mc1_dis_ufm     : in     vl_logic;
        mc1_done_phase  : in     vl_logic_vector(1 downto 0);
        mc1_dsr_fctrl   : in     vl_logic_vector(1 downto 0);
        mc1_en_cfgstdby : in     vl_logic;
        mc1_en_cibstdby : in     vl_logic;
        mc1_en_cibwake  : in     vl_logic;
        mc1_en_i2cwake  : in     vl_logic;
        mc1_ents        : in     vl_logic;
        mc1_er1_exist   : in     vl_logic;
        mc1_er2_exist   : in     vl_logic;
        mc1_goe         : in     vl_logic;
        mc1_goe_phase   : in     vl_logic_vector(1 downto 0);
        mc1_gsr_phase   : in     vl_logic_vector(1 downto 0);
        mc1_gsrn        : in     vl_logic;
        mc1_gsrn_cib    : in     vl_logic;
        mc1_gsrn_inv    : in     vl_logic;
        mc1_gsrn_sync   : in     vl_logic;
        mc1_gwe         : in     vl_logic;
        mc1_gwe_phase   : in     vl_logic_vector(1 downto 0);
        mc1_i2c_persist : in     vl_logic;
        mc1_mclk_cib    : in     vl_logic_vector(6 downto 0);
        mc1_mib         : in     vl_logic;
        mc1_mspi_addr   : in     vl_logic_vector(7 downto 0);
        mc1_mspi_persist: in     vl_logic;
        mc1_mspi_sedaddr: in     vl_logic_vector(15 downto 0);
        mc1_pll_set     : in     vl_logic;
        mc1_ppt_qout    : in     vl_logic_vector(7 downto 0);
        mc1_sed_once    : in     vl_logic;
        mc1_sed_always  : in     vl_logic;
        mc1_sed_clk     : in     vl_logic_vector(6 downto 0);
        mc1_sed_en      : in     vl_logic_vector(1 downto 0);
        mc1_source_sel  : in     vl_logic;
        mc1_sspi_persist: in     vl_logic;
        mc1_stdby_bg    : in     vl_logic_vector(1 downto 0);
        mc1_syn_ext_done: in     vl_logic;
        mc1_syn_src     : in     vl_logic;
        mc1_tsinv       : in     vl_logic;
        mc1_user_timer  : in     vl_logic;
        mc1_wl_slew     : in     vl_logic;
        cib_i2c_scl_i   : in     vl_logic;
        cib_i2c_sda_i   : in     vl_logic;
        cib_sspi_csn    : in     vl_logic;
        jtdo            : in     vl_logic_vector(2 downto 1);
        cib_auto_reboot : in     vl_logic;
        cib_clr_flag    : in     vl_logic;
        cib_mspi_addr   : in     vl_logic_vector(7 downto 0);
        cib_osc_dis     : in     vl_logic;
        cib_stdby       : in     vl_logic;
        cib_stdby_clk   : in     vl_logic;
        cib_timeout     : in     vl_logic;
        cib_ts_all      : in     vl_logic;
        gsrn_sync_clk   : in     vl_logic;
        pll_lock        : in     vl_logic;
        sed_clk         : in     vl_logic;
        sed_enable      : in     vl_logic;
        sed_frcerr      : in     vl_logic;
        sed_mode        : in     vl_logic;
        sed_start       : in     vl_logic;
        user_clk        : in     vl_logic;
        usr_gsr         : in     vl_logic;
        es_i            : in     vl_logic_vector(8 downto 0);
        fl_c_bl         : in     vl_logic_vector(3 downto 0);
        fl_dout         : in     vl_logic_vector(63 downto 0);
        fl_lastcol      : in     vl_logic_vector(3 downto 0);
        fl_neg_edge_det : in     vl_logic;
        fl_ready_vfy    : in     vl_logic;
        fl_vwlp_active  : in     vl_logic;
        fl_well_active  : in     vl_logic;
        fl_ready        : in     vl_logic;
        fl_l_row_cfg    : in     vl_logic;
        fl_l_row_ufm    : in     vl_logic;
        scan2_out       : in     vl_logic;
        scanen          : in     vl_logic;
        i2cbr_1st       : in     vl_logic_vector(9 downto 0);
        i2cbr_2nd       : in     vl_logic_vector(9 downto 0);
        i2ccmdr_1st     : in     vl_logic_vector(7 downto 2);
        i2ccmdr_2nd     : in     vl_logic_vector(7 downto 2);
        i2ccr1_1st      : in     vl_logic_vector(7 downto 2);
        i2ccr1_2nd      : in     vl_logic_vector(7 downto 2);
        i2ctxdr_1st     : in     vl_logic_vector(7 downto 0);
        i2ctxdr_2nd     : in     vl_logic_vector(7 downto 0);
        spibr           : in     vl_logic_vector(5 downto 0);
        spicr0          : in     vl_logic_vector(7 downto 0);
        spicr1          : in     vl_logic_vector(7 downto 4);
        spicr2          : in     vl_logic_vector(7 downto 0);
        spicsr          : in     vl_logic_vector(7 downto 0);
        spitxdr         : in     vl_logic_vector(7 downto 0);
        wbccr           : in     vl_logic_vector(7 downto 6);
        wbctxdr         : in     vl_logic_vector(7 downto 0);
        stb_i2cbr_1st   : in     vl_logic;
        stb_i2cbr_2nd   : in     vl_logic;
        stb_i2ccmdr_1st : in     vl_logic;
        stb_i2ccmdr_2nd : in     vl_logic;
        stb_i2ccr1_1st  : in     vl_logic;
        stb_i2ccr1_2nd  : in     vl_logic;
        stb_i2cgcdr_1st : in     vl_logic;
        stb_i2cgcdr_2nd : in     vl_logic;
        stb_i2crxdr_1st : in     vl_logic;
        stb_i2crxdr_2nd : in     vl_logic;
        stb_i2ctxdr_1st : in     vl_logic;
        stb_i2ctxdr_2nd : in     vl_logic;
        stb_spibr       : in     vl_logic;
        stb_spicr0      : in     vl_logic;
        stb_spicr1      : in     vl_logic;
        stb_spicr2      : in     vl_logic;
        stb_spicsr      : in     vl_logic;
        stb_spirxdr     : in     vl_logic;
        stb_spitxdr     : in     vl_logic;
        stb_wbccr       : in     vl_logic;
        stb_wbcrxdr     : in     vl_logic;
        stb_wbctxdr     : in     vl_logic;
        sciclk_tree     : in     vl_logic;
        sciclk          : in     vl_logic
    );
end config_plus;
