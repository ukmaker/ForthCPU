library verilog;
use verilog.vl_types.all;
entity SEH_OR2_2 is
    port(
        X               : out    vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic
    );
end SEH_OR2_2;
