library verilog;
use verilog.vl_types.all;
entity vlov1s is
    port(
        Z               : out    vl_logic
    );
end vlov1s;
