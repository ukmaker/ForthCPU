library verilog;
use verilog.vl_types.all;
entity DNEQ_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end DNEQ_UDP;
