library verilog;
use verilog.vl_types.all;
entity TGM4_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end TGM4_UDP;
