library verilog;
use verilog.vl_types.all;
entity memctrl is
    port(
        erasprgmtmr_test: out    vl_logic;
        wrrdvid1_iflg   : out    vl_logic;
        wrrdvid2_iflg   : out    vl_logic;
        wrrdvid3_iflg   : out    vl_logic;
        wrrdvid4_iflg   : out    vl_logic;
        wrrdvid5_iflg   : out    vl_logic;
        wrrdvid6_iflg   : out    vl_logic;
        wrrdvid7_iflg   : out    vl_logic;
        wrrdvid8_iflg   : out    vl_logic;
        vidbyte1_sel    : out    vl_logic;
        mfg_load_addrlat: out    vl_logic;
        mfg_load_datareg: out    vl_logic;
        readmfg_drvmcbus: out    vl_logic;
        cfgtrim_load_addrlat: out    vl_logic;
        cfgtrim_load_datareg: out    vl_logic;
        cfgtrim_drvmcbus: out    vl_logic;
        cfgarray_data_enable: out    vl_logic;
        cfgtrim_sel_datareg: out    vl_logic;
        cfg_load_shdwregaddrlat: out    vl_logic;
        cfgshdw_ld_m_latch: out    vl_logic;
        cfgshdw_ld_m_latch_iawp: out    vl_logic;
        cfgshdw_ld_s_latch: out    vl_logic;
        nscb_cfgmshdw_drvmcbus: out    vl_logic;
        mc_twifl_data   : out    vl_logic_vector(7 downto 0);
        faultlog_sel_3wi: out    vl_logic;
        flut_col_addr   : out    vl_logic_vector(2 downto 0);
        flut_row_addr   : out    vl_logic_vector(3 downto 0);
        flut_load_datareg: out    vl_logic;
        faultlog_load_soft_datareg: out    vl_logic;
        flut_drvmcbus   : out    vl_logic;
        faultlog_in_progress: out    vl_logic;
        faultlog_full   : out    vl_logic;
        eep_shdw_ready  : out    vl_logic;
        i2csa_load_datareg: out    vl_logic;
        i2csa_drvmcbus  : out    vl_logic;
        readid_drvmcbus : out    vl_logic;
        done_sel_array  : out    vl_logic;
        i2csa_sel_array : out    vl_logic;
        cfg_sel_array   : out    vl_logic;
        flut_sel_array  : out    vl_logic;
        trim_sel_array  : out    vl_logic;
        enable_prgrm    : out    vl_logic;
        enable_erase    : out    vl_logic;
        enable_dischrg  : out    vl_logic;
        enable_verify   : out    vl_logic;
        noack           : out    vl_logic;
        safestate       : out    vl_logic;
        tristpad_iflg   : out    vl_logic;
        en_i2c_dat      : out    vl_logic;
        mc_mcb_out      : out    vl_logic_vector(7 downto 0);
        mc_drvmcbus     : out    vl_logic;
        measctrl_load_addrlat: out    vl_logic;
        measctrl_load_datalat: out    vl_logic;
        measresult_drvmcbus: out    vl_logic;
        ctrl_vhien      : out    vl_logic;
        trim_load_shdwregaddrlat: out    vl_logic;
        trimshdw_ld_latch: out    vl_logic;
        trimshdw_drvmcbus: out    vl_logic;
        north_keeper_drvmcbus: out    vl_logic;
        reset_in_b      : in     vl_logic;
        clk_8mhz        : in     vl_logic;
        testentimer     : in     vl_logic;
        testclken       : in     vl_logic;
        mc_mcb_in       : in     vl_logic_vector(7 downto 0);
        wrir_in         : in     vl_logic;
        wrd_in          : in     vl_logic;
        rdd_in          : in     vl_logic;
        donebit         : in     vl_logic;
        i2csadone       : in     vl_logic;
        mfg_mode        : in     vl_logic;
        gpiopincfgwrprotec_b: in     vl_logic;
        twi_start       : in     vl_logic;
        twi_wdat_write_reg: in     vl_logic;
        twi_rdat_read   : in     vl_logic;
        twi_rdat_data_from_latch: in     vl_logic_vector(7 downto 0);
        twi_flid_shdw   : in     vl_logic_vector(7 downto 0);
        twi_fl_record   : in     vl_logic;
        twi_fl_soft     : in     vl_logic;
        erase_slot      : in     vl_logic_vector(3 downto 0);
        erase_range     : in     vl_logic_vector(1 downto 0);
        progm_slot      : in     vl_logic_vector(3 downto 0);
        progm_range     : in     vl_logic_vector(1 downto 0);
        fl_prgm_slot    : in     vl_logic_vector(3 downto 0);
        fl_prgm_range   : in     vl_logic_vector(1 downto 0);
        fsafe           : in     vl_logic
    );
end memctrl;
