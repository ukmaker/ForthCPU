library verilog;
use verilog.vl_types.all;
entity pcs_dual_dp is
    port(
        bus8bit_sel     : in     vl_logic;
        bist_rx_data_sel: in     vl_logic;
        char_test_mode  : in     vl_logic;
        char_test_data  : in     vl_logic_vector(9 downto 0);
        ebrd_clk        : in     vl_logic_vector(1 downto 0);
        fbw_clk         : in     vl_logic_vector(1 downto 0);
        ff_tx_d_0       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_1       : in     vl_logic_vector(23 downto 0);
        ffc_ei_en       : in     vl_logic_vector(1 downto 0);
        ffc_enable_cgalign: in     vl_logic_vector(1 downto 0);
        ffc_fb_loopback : in     vl_logic_vector(1 downto 0);
        ffc_pcie_det_en : in     vl_logic_vector(1 downto 0);
        ffc_pcie_ct     : in     vl_logic_vector(1 downto 0);
        pfifow_clr      : in     vl_logic_vector(1 downto 0);
        pfifor_clr      : in     vl_logic_vector(1 downto 0);
        pfifo_clr_sel   : in     vl_logic;
        ffc_rxpwdnb     : in     vl_logic_vector(1 downto 0);
        ffc_sb_inv_rx   : in     vl_logic_vector(1 downto 0);
        ffc_sb_pfifo_lp : in     vl_logic_vector(1 downto 0);
        ffc_signal_detect: in     vl_logic_vector(1 downto 0);
        ffc_txpwdnb     : in     vl_logic_vector(1 downto 0);
        ffc_rx_div11_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_div11_mode: in     vl_logic_vector(1 downto 0);
        ffc_rx_rate_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_rate_mode: in     vl_logic_vector(1 downto 0);
        ffc_rx_gear_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_gear_mode: in     vl_logic_vector(1 downto 0);
        ffc_cdr_en_bitslip: in     vl_logic_vector(1 downto 0);
        fmbist_data     : in     vl_logic_vector(9 downto 0);
        bist_ch_sel     : in     vl_logic;
        force_int       : in     vl_logic;
        rxf_clk         : in     vl_logic_vector(1 downto 0);
        txf_clk         : in     vl_logic_vector(1 downto 0);
        ffc_ldr_core2tx_en: in     vl_logic_vector(1 downto 0);
        mc1_chif_ctl_ch0: in     vl_logic_vector(263 downto 0);
        mc1_chif_ctl_ch1: in     vl_logic_vector(263 downto 0);
        mc1_ser_ctl_ch0 : in     vl_logic_vector(87 downto 0);
        mc1_ser_ctl_ch1 : in     vl_logic_vector(87 downto 0);
        pci_connect     : in     vl_logic_vector(1 downto 0);
        pcs_ctl_3_dl_02 : in     vl_logic_vector(7 downto 0);
        plol            : in     vl_logic;
        rlol            : in     vl_logic_vector(1 downto 0);
        rlos            : in     vl_logic_vector(1 downto 0);
        pci_det_done    : in     vl_logic_vector(1 downto 0);
        rxr_clk         : in     vl_logic_vector(1 downto 0);
        rx_d_sd_0       : in     vl_logic_vector(9 downto 0);
        rx_d_sd_1       : in     vl_logic_vector(9 downto 0);
        sciaddr         : in     vl_logic_vector(5 downto 0);
        sciwdata        : in     vl_logic_vector(7 downto 0);
        scird           : in     vl_logic;
        cyawstn         : in     vl_logic;
        sciench0        : in     vl_logic;
        sciench1        : in     vl_logic;
        sciselch0       : in     vl_logic;
        sciselch1       : in     vl_logic;
        ser_sts_2_ch_27_0: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_1: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_0: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_1: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_0: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_1: in     vl_logic_vector(7 downto 0);
        txp_clk         : in     vl_logic_vector(1 downto 0);
        xge_mode        : in     vl_logic;
        done_cfg        : in     vl_logic;
        reg_load        : in     vl_logic;
        goe_r2          : in     vl_logic;
        goe_load        : in     vl_logic;
        rstb_txf        : in     vl_logic_vector(1 downto 0);
        rstb_txp        : in     vl_logic_vector(1 downto 0);
        rstb_ebrd       : in     vl_logic_vector(1 downto 0);
        rstb_rxr        : in     vl_logic_vector(1 downto 0);
        rstb_fbw        : in     vl_logic_vector(1 downto 0);
        rstb_rxf        : in     vl_logic_vector(1 downto 0);
        ff_rx_d_0       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_1       : out    vl_logic_vector(23 downto 0);
        pci_det_en      : out    vl_logic_vector(1 downto 0);
        ffs_cc_overrun  : out    vl_logic_vector(1 downto 0);
        ffs_cc_underrun : out    vl_logic_vector(1 downto 0);
        ffs_ls_sync_status: out    vl_logic_vector(1 downto 0);
        ffs_rxfbfifo_error: out    vl_logic_vector(1 downto 0);
        ffs_txfbfifo_error: out    vl_logic_vector(1 downto 0);
        ffs_rlos        : out    vl_logic_vector(1 downto 0);
        ffs_pcie_done   : out    vl_logic_vector(1 downto 0);
        ffs_pcie_con    : out    vl_logic_vector(1 downto 0);
        pcie_mode       : out    vl_logic_vector(1 downto 0);
        pcie_phystatus  : out    vl_logic_vector(1 downto 0);
        pcie_rxvalid    : out    vl_logic_vector(1 downto 0);
        skp_added       : out    vl_logic_vector(1 downto 0);
        skp_deleted     : out    vl_logic_vector(1 downto 0);
        full_d          : out    vl_logic_vector(1 downto 0);
        empty_d         : out    vl_logic_vector(1 downto 0);
        rx_ch           : out    vl_logic_vector(1 downto 0);
        tx_d_sd_0       : out    vl_logic_vector(9 downto 0);
        tx_d_sd_1       : out    vl_logic_vector(9 downto 0);
        sciint_10       : out    vl_logic_vector(1 downto 0);
        scirdata_01     : out    vl_logic_vector(7 downto 0);
        rst_ctl_1_ch_1f_0: out    vl_logic_vector(7 downto 0);
        rst_ctl_1_ch_1f_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_8_ch_17_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_8_ch_17_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_9_ch_18_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_9_ch_18_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_10_ch_19_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_10_ch_19_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_11_ch_1a_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_11_ch_1a_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_12_ch_1b_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_12_ch_1b_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_13_ch_1c_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_13_ch_1c_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_14_ch_1d_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_14_ch_1d_1: out    vl_logic_vector(7 downto 0);
        pcs_ctl_3_ch_02_710: out    vl_logic_vector(3 downto 0);
        pcs_ctl_3_ch_02_32: out    vl_logic_vector(3 downto 0);
        tobist_data     : out    vl_logic_vector(9 downto 0);
        pci_det_ct      : out    vl_logic_vector(1 downto 0);
        pci_ei_en       : out    vl_logic_vector(1 downto 0);
        cdr_en_bitslip0 : out    vl_logic;
        cdr_en_bitslip1 : out    vl_logic;
        cout            : out    vl_logic_vector(15 downto 0);
        ser_mem_ch0     : out    vl_logic_vector(87 downto 0);
        ser_mem_ch1     : out    vl_logic_vector(87 downto 0)
    );
end pcs_dual_dp;
