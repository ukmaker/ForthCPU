library verilog;
use verilog.vl_types.all;
entity config_core is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 0;
        DECRYPTION      : integer := 0
    );
    port(
        done_gwe        : out    vl_logic;
        gsrn_sync       : out    vl_logic;
        gsrn            : out    vl_logic;
        goe             : out    vl_logic;
        en_pupn         : out    vl_logic;
        freeze_io       : out    vl_logic;
        freeze_mib      : out    vl_logic;
        pcs_rstn        : out    vl_logic;
        jtck            : out    vl_logic;
        int_spi_mclk    : out    vl_logic;
        int_spi_data    : out    vl_logic_vector(15 downto 0);
        int_spi_mcsn    : out    vl_logic_vector(7 downto 0);
        tlreset         : out    vl_logic;
        bsrclk          : out    vl_logic;
        shiftdr_bs      : out    vl_logic;
        updatedr_bs     : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        ac_mode         : out    vl_logic;
        ac_clear        : out    vl_logic;
        ac_test         : out    vl_logic;
        tdi_bscan       : out    vl_logic;
        ts_all          : out    vl_logic;
        jtag_persist    : out    vl_logic;
        progn_persist   : out    vl_logic;
        initn_persist   : out    vl_logic;
        donep_persist   : out    vl_logic;
        sram_asr_clk    : out    vl_logic;
        sram_asr_in     : out    vl_logic;
        sram_asr_rst    : out    vl_logic;
        sram_asr_en_incr: out    vl_logic;
        sram_asr_shift_1st: out    vl_logic;
        sram_asr_shift_2nd: out    vl_logic;
        sram_asr_shift_3rd: out    vl_logic;
        sf_ppt_addr     : out    vl_logic_vector(3 downto 0);
        sram_wl_str     : out    vl_logic;
        sram_data_wr    : out    vl_logic;
        cfg_addr_slew   : out    vl_logic;
        cfg_data_cap    : out    vl_logic;
        cfg_data_flt    : out    vl_logic;
        cfg_data_pre    : out    vl_logic;
        dsr_clk         : out    vl_logic;
        dsr_din         : out    vl_logic_vector(63 downto 0);
        dsr_upd_lat     : out    vl_logic;
        dsr_cap         : out    vl_logic;
        dsr_rst_n       : out    vl_logic;
        dsr_shift       : out    vl_logic_vector(1 downto 0);
        ef_en           : out    vl_logic;
        ef_rw           : out    vl_logic;
        ef_execute      : out    vl_logic;
        ef_row_addr     : out    vl_logic_vector(4 downto 0);
        ef_col_addr     : out    vl_logic_vector(6 downto 0);
        mfg_ef_margin   : out    vl_logic;
        mfg_ef_atest    : out    vl_logic_vector(1 downto 0);
        trim_ef_acntl   : out    vl_logic_vector(7 downto 0);
        instr_dts       : out    vl_logic;
        start_dts       : out    vl_logic;
        dtsclk          : out    vl_logic;
        initn_o         : out    vl_logic;
        initn_oe        : out    vl_logic;
        donep_o         : out    vl_logic;
        donep_oe        : out    vl_logic;
        mcsn_o          : out    vl_logic_vector(7 downto 0);
        mcsn_oe         : out    vl_logic_vector(7 downto 0);
        mclk_o          : out    vl_logic;
        mclk_oe         : out    vl_logic;
        sspi_so         : out    vl_logic;
        sspi_oe         : out    vl_logic;
        mclk_byp_o      : out    vl_logic;
        mclk_byp_oe     : out    vl_logic;
        data_o          : out    vl_logic_vector(15 downto 0);
        data_oe         : out    vl_logic_vector(15 downto 0);
        docson_o        : out    vl_logic;
        docson_oe       : out    vl_logic;
        busy_o          : out    vl_logic;
        busy_oe         : out    vl_logic;
        tdo_o           : out    vl_logic;
        tdo_oe          : out    vl_logic;
        sda_out_pad     : out    vl_logic;
        sda_oe_pad      : out    vl_logic;
        scl_out_pad     : out    vl_logic;
        scl_oe_pad      : out    vl_logic;
        isptcy_ener1    : out    vl_logic;
        isptcy_ener2    : out    vl_logic;
        isptcy_resetb   : out    vl_logic;
        isptcy_shcap    : out    vl_logic;
        isptcy_update   : out    vl_logic;
        isptcy_rtier1   : out    vl_logic;
        isptcy_rtier2   : out    vl_logic;
        isptcy_tdi      : out    vl_logic;
        sed_auto_done_cib: out    vl_logic;
        sed_clk_cib     : out    vl_logic;
        sed_done_cib    : out    vl_logic;
        sed_busy_cib    : out    vl_logic;
        sed_err_cib     : out    vl_logic;
        cfg_done_cib    : out    vl_logic;
        freeze_io_cib   : out    vl_logic;
        last_addr_cib   : out    vl_logic_vector(15 downto 0);
        persist_out_cib : out    vl_logic_vector(15 downto 0);
        usrclk_cib      : out    vl_logic;
        sda_out_cib     : out    vl_logic;
        sda_oe_cib      : out    vl_logic;
        scl_out_cib     : out    vl_logic;
        scl_oe_cib      : out    vl_logic;
        mcsn_o_cib      : out    vl_logic_vector(7 downto 0);
        mcsn_oe_cib     : out    vl_logic_vector(7 downto 0);
        mclk_o_2nd      : out    vl_logic;
        mclk_oe_2nd     : out    vl_logic;
        mosi_o_2nd      : out    vl_logic;
        mosi_oe_2nd     : out    vl_logic;
        miso_o_2nd      : out    vl_logic;
        miso_oe_2nd     : out    vl_logic;
        es_o            : out    vl_logic_vector(35 downto 0);
        pcs_o           : out    vl_logic_vector(27 downto 0);
        iscan_en        : out    vl_logic_vector(7 downto 0);
        i2crxdr_1st     : out    vl_logic_vector(7 downto 0);
        i2cgcdr_1st     : out    vl_logic_vector(7 downto 0);
        i2csr_1st       : out    vl_logic_vector(7 downto 0);
        i2c_wkup_1st    : out    vl_logic;
        i2crxdr_2nd     : out    vl_logic_vector(7 downto 0);
        i2cgcdr_2nd     : out    vl_logic_vector(7 downto 0);
        i2csr_2nd       : out    vl_logic_vector(7 downto 0);
        i2c_wkup_2nd    : out    vl_logic;
        wbcsr           : out    vl_logic_vector(7 downto 0);
        wbcrxdr         : out    vl_logic_vector(7 downto 0);
        spisr           : out    vl_logic_vector(7 downto 0);
        spirxdr         : out    vl_logic_vector(7 downto 0);
        spi_wkup        : out    vl_logic;
        stdby_ena       : out    vl_logic;
        dev_stdby_exec  : out    vl_logic;
        dev_sleep_exec  : out    vl_logic;
        dev_wkup_exec   : out    vl_logic;
        ppt_en          : out    vl_logic;
        ppt_rowsel      : out    vl_logic;
        ppt_pset        : out    vl_logic;
        row             : out    vl_logic_vector(14 downto 0);
        ufm_row_sel_all : out    vl_logic;
        ufm_row_sel_none: out    vl_logic;
        cfg_row_sel_all : out    vl_logic;
        cfg_row_sel_none: out    vl_logic;
        trim_row_sel_all: out    vl_logic;
        trim_row_sel_none: out    vl_logic;
        feat_row_sel_all: out    vl_logic;
        feat_row_sel_none: out    vl_logic;
        era_ufm         : out    vl_logic;
        era_cfg         : out    vl_logic;
        era_trim        : out    vl_logic;
        era_feat        : out    vl_logic;
        prg_ufm         : out    vl_logic;
        prg_cfg         : out    vl_logic;
        prg_tf          : out    vl_logic;
        read_ufm        : out    vl_logic;
        read_cfg        : out    vl_logic;
        read_tf         : out    vl_logic;
        erase_setup     : out    vl_logic;
        erapdis         : out    vl_logic;
        erase_pulse     : out    vl_logic;
        pwtc_well       : out    vl_logic;
        prg_pulse       : out    vl_logic_vector(3 downto 0);
        prog_disch      : out    vl_logic;
        prg_pwtc        : out    vl_logic;
        en_vreg_mon     : out    vl_logic;
        era_ver         : out    vl_logic;
        scp             : out    vl_logic;
        softprg         : out    vl_logic;
        verify          : out    vl_logic;
        flash_en        : out    vl_logic;
        reg_enable      : out    vl_logic;
        scpv            : out    vl_logic;
        subrow_mvena_ufm: out    vl_logic;
        subrow_mvenall_ufm: out    vl_logic;
        subrow_hvena_ufm: out    vl_logic;
        subrow_hvenall_ufm: out    vl_logic;
        subrow_mvena_cfg: out    vl_logic;
        subrow_mvenall_cfg: out    vl_logic;
        subrow_hvena_cfg: out    vl_logic;
        subrow_hvenall_cfg: out    vl_logic;
        subrow_mvena_tf : out    vl_logic;
        subrow_hvena_tf : out    vl_logic;
        sa_enall        : out    vl_logic;
        sa_ena          : out    vl_logic;
        prgdrv_enall    : out    vl_logic;
        prgdrv_ena      : out    vl_logic;
        col_shift       : out    vl_logic;
        col_rst         : out    vl_logic;
        colstart        : out    vl_logic_vector(3 downto 0);
        readpart        : out    vl_logic_vector(3 downto 0);
        wor_eval        : out    vl_logic;
        wand_eval       : out    vl_logic;
        capture_dout    : out    vl_logic;
        src_clamp       : out    vl_logic;
        drain_ctrl      : out    vl_logic;
        sel_6p5v        : out    vl_logic;
        prestep_in_neg  : out    vl_logic_vector(2 downto 0);
        step_in_neg     : out    vl_logic_vector(2 downto 0);
        fl_ready_rst    : out    vl_logic;
        mfg_margin_en   : out    vl_logic;
        flash_clk_mfg   : out    vl_logic;
        mux32_out1      : out    vl_logic;
        mux32_out2      : out    vl_logic;
        trim_osc        : out    vl_logic_vector(7 downto 0);
        trim_bg         : out    vl_logic_vector(15 downto 0);
        trim_spare      : out    vl_logic_vector(63 downto 0);
        mfg_pll_out     : out    vl_logic_vector(1 downto 0);
        mfg_spare       : out    vl_logic_vector(47 downto 0);
        por             : in     vl_logic;
        intclk          : in     vl_logic;
        sleep_mode      : in     vl_logic;
        CHIPID          : in     vl_logic_vector(7 downto 0);
        CTRL0_DEFAULT   : in     vl_logic_vector(31 downto 0);
        CRC32_DEFAULT   : in     vl_logic_vector(31 downto 0);
        UCODE_DEFAULT   : in     vl_logic_vector(31 downto 0);
        NDUM_DEFAULT    : in     vl_logic_vector(3 downto 0);
        ASSP_EN         : in     vl_logic;
        HFC_EN          : in     vl_logic;
        ENC_ONLY_EN     : in     vl_logic;
        IDCODE0         : in     vl_logic_vector(31 downto 0);
        ASR_LENGTH      : in     vl_logic_vector(13 downto 0);
        DSR_LENGTH      : in     vl_logic_vector(15 downto 0);
        EBR_ROW         : in     vl_logic_vector(3 downto 0);
        PLC_COL         : in     vl_logic_vector(9 downto 0);
        RES_COL         : in     vl_logic_vector(2 downto 0);
        RES_COL_NUM     : in     vl_logic_vector(39 downto 0);
        INT_SPI_CTRL    : in     vl_logic_vector(1 downto 0);
        fsafe           : in     vl_logic;
        scanen          : in     vl_logic;
        int_spi_din     : in     vl_logic_vector(15 downto 0);
        bscan_out       : in     vl_logic;
        asr_rmr_out     : in     vl_logic;
        dsr_rcr_out     : in     vl_logic_vector(7 downto 0);
        iscan_out       : in     vl_logic_vector(7 downto 0);
        hfc_select_pin  : in     vl_logic;
        cclk_pin        : in     vl_logic;
        mclk_pin        : in     vl_logic;
        gsrn_pin        : in     vl_logic;
        cs0n            : in     vl_logic;
        cs1n            : in     vl_logic;
        din             : in     vl_logic_vector(15 downto 0);
        di              : in     vl_logic;
        done_pin        : in     vl_logic;
        initn_pin       : in     vl_logic;
        cfg_pin         : in     vl_logic_vector(2 downto 0);
        programn_pin    : in     vl_logic;
        writen_pin      : in     vl_logic;
        tck_pin         : in     vl_logic;
        tdi_pin         : in     vl_logic;
        tms_pin         : in     vl_logic;
        jtagenb_pin     : in     vl_logic;
        sda_in_pad      : in     vl_logic;
        scl_in_pad      : in     vl_logic;
        pwr_save_mode   : in     vl_logic;
        mc1_sed_auto_rboot: in     vl_logic;
        mc1_sed_enable  : in     vl_logic_vector(1 downto 0);
        mc1_sed_clk     : in     vl_logic_vector(6 downto 0);
        mc1_sed_always  : in     vl_logic;
        mc1_sed_sleep   : in     vl_logic;
        mc1_sed_once    : in     vl_logic;
        mc1_dsr_fctrl   : in     vl_logic_vector(1 downto 0);
        mc1_done_phase  : in     vl_logic_vector(3 downto 0);
        mc1_goe_phase   : in     vl_logic_vector(2 downto 0);
        mc1_gsr_phase   : in     vl_logic_vector(2 downto 0);
        mc1_gwe_phase   : in     vl_logic_vector(2 downto 0);
        mc1_gsrn        : in     vl_logic;
        mc1_gsrn_inv    : in     vl_logic;
        mc1_gsrn_sync   : in     vl_logic;
        mc1_gwe         : in     vl_logic;
        mc1_sync_ext_done: in     vl_logic;
        mc1_sync_source : in     vl_logic;
        mc1_goe         : in     vl_logic;
        mc1_mib         : in     vl_logic;
        mc1_pcs         : in     vl_logic;
        mc1_persist_cap : in     vl_logic;
        mc1_pll_chk     : in     vl_logic_vector(7 downto 0);
        mc1_pupn        : in     vl_logic;
        mc1_user_gsrn   : in     vl_logic;
        mc1_source_sel  : in     vl_logic;
        mc1_mspi_addr   : in     vl_logic_vector(15 downto 0);
        mc1_mspi_sed_addr: in     vl_logic_vector(15 downto 0);
        mc1_en_tsall    : in     vl_logic;
        mc1_tsall_inv   : in     vl_logic;
        mc1_usr_clk     : in     vl_logic_vector(6 downto 0);
        mc1_er1_exist   : in     vl_logic;
        mc1_er2_exist   : in     vl_logic;
        mc1_dts_clk     : in     vl_logic;
        mc1_sleep_gsrn  : in     vl_logic;
        mc1_sleep_gwe   : in     vl_logic;
        mc1_sleep_pupn  : in     vl_logic;
        mc1_sleep_fio   : in     vl_logic;
        mc1_persist_mspi: in     vl_logic;
        mc1_persist_sspi: in     vl_logic;
        mc1_persist_i2c : in     vl_logic;
        mc1_persist_cpu8: in     vl_logic;
        mc1_persist_cpu16: in     vl_logic;
        mc1_bl_float    : in     vl_logic;
        mc1_wl_slew     : in     vl_logic;
        mc1_ppt_bits    : in     vl_logic_vector(7 downto 0);
        isptracy_er1_out: in     vl_logic;
        isptracy_er2_out: in     vl_logic;
        cib_auto_reboot : in     vl_logic;
        cib_mspim_addr  : in     vl_logic_vector(15 downto 0);
        cib_tsall       : in     vl_logic;
        cib_persist_in  : in     vl_logic_vector(15 downto 0);
        cib_pll_lock    : in     vl_logic_vector(7 downto 0);
        cib_sed_clk     : in     vl_logic;
        cib_sed_en      : in     vl_logic;
        cib_sed_frcerr  : in     vl_logic;
        cib_sed_mode    : in     vl_logic;
        cib_sed_start   : in     vl_logic;
        cib_wkup_clk    : in     vl_logic;
        cib_user_gsr    : in     vl_logic;
        cib_mcsn_sel    : in     vl_logic;
        sda_in_cib      : in     vl_logic;
        scl_in_cib      : in     vl_logic;
        sclk_i_2nd      : in     vl_logic;
        mosi_i_2nd      : in     vl_logic;
        miso_i_2nd      : in     vl_logic;
        scsn_2nd_cib    : in     vl_logic;
        bg_cmp_out      : in     vl_logic;
        bg_rdy          : in     vl_logic;
        proc_ring_osc   : in     vl_logic;
        dts_out         : in     vl_logic_vector(31 downto 0);
        es_i            : in     vl_logic_vector(8 downto 0);
        pcs_i           : in     vl_logic_vector(7 downto 0);
        pcs_stat        : in     vl_logic_vector(2 downto 0);
        device          : in     vl_logic_vector(2 downto 0);
        c_bl            : in     vl_logic_vector(3 downto 0);
        fl_dout         : in     vl_logic_vector(63 downto 0);
        lastcol         : in     vl_logic_vector(3 downto 0);
        fl_ready        : in     vl_logic;
        l_row_cfg       : in     vl_logic;
        l_row_ufm       : in     vl_logic;
        neg_edge_det    : in     vl_logic;
        vwlp_active     : in     vl_logic;
        ready_vfy       : in     vl_logic;
        well_active     : in     vl_logic;
        ef_do           : in     vl_logic;
        sf_asr_out      : in     vl_logic;
        wb_clk_i        : in     vl_logic;
        wb_clk_nt       : in     vl_logic;
        spicr0          : in     vl_logic_vector(7 downto 0);
        spicr1          : in     vl_logic_vector(7 downto 0);
        spicr2          : in     vl_logic_vector(7 downto 0);
        spibr           : in     vl_logic_vector(7 downto 0);
        spicsr          : in     vl_logic_vector(7 downto 0);
        spitxdr         : in     vl_logic_vector(7 downto 0);
        wb_spicr0_wt    : in     vl_logic;
        wb_spicr1_wt    : in     vl_logic;
        wb_spicr2_wt    : in     vl_logic;
        wb_spibr_wt     : in     vl_logic;
        wb_spicsr_wt    : in     vl_logic;
        wb_spitxdr_wt   : in     vl_logic;
        wb_spirxdr_rd   : in     vl_logic;
        wbccr1          : in     vl_logic_vector(7 downto 0);
        wbctxdr         : in     vl_logic_vector(7 downto 0);
        wb_wbccr1_wt    : in     vl_logic;
        wb_wbctxdr_wt   : in     vl_logic;
        wb_wbcrxdr_rd   : in     vl_logic;
        i2ccr1_1st      : in     vl_logic_vector(7 downto 0);
        i2ccmdr_1st     : in     vl_logic_vector(7 downto 0);
        i2ctxdr_1st     : in     vl_logic_vector(7 downto 0);
        i2cbr_1st       : in     vl_logic_vector(9 downto 0);
        wb_i2ccr1_wt_1st: in     vl_logic;
        wb_i2ccmdr_wt_1st: in     vl_logic;
        wb_i2cbr_wt_1st : in     vl_logic;
        wb_i2ctxdr_wt_1st: in     vl_logic;
        wb_i2crxdr_rd_1st: in     vl_logic;
        wb_i2cgcdr_rd_1st: in     vl_logic;
        i2ccr1_2nd      : in     vl_logic_vector(7 downto 0);
        i2ccmdr_2nd     : in     vl_logic_vector(7 downto 0);
        i2ctxdr_2nd     : in     vl_logic_vector(7 downto 0);
        i2cbr_2nd       : in     vl_logic_vector(9 downto 0);
        wb_i2ccr1_wt_2nd: in     vl_logic;
        wb_i2ccmdr_wt_2nd: in     vl_logic;
        wb_i2cbr_wt_2nd : in     vl_logic;
        wb_i2ctxdr_wt_2nd: in     vl_logic;
        wb_i2crxdr_rd_2nd: in     vl_logic;
        wb_i2cgcdr_rd_2nd: in     vl_logic
    );
end config_core;
