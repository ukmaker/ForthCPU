library verilog;
use verilog.vl_types.all;
entity pcs_dual is
    port(
        cin             : in     vl_logic_vector(11 downto 0);
        cyawstn         : in     vl_logic;
        ff_ebrd_clk     : in     vl_logic_vector(1 downto 0);
        ff_rxi_clk      : in     vl_logic_vector(1 downto 0);
        ff_tx_d_0       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_1       : in     vl_logic_vector(23 downto 0);
        ff_txi_clk      : in     vl_logic_vector(1 downto 0);
        ffc_ei_en       : in     vl_logic_vector(1 downto 0);
        ffc_enable_cgalign: in     vl_logic_vector(1 downto 0);
        ffc_fb_loopback : in     vl_logic_vector(1 downto 0);
        ffc_rx_lane_rst : in     vl_logic_vector(1 downto 0);
        ffc_tx_lane_rst : in     vl_logic_vector(1 downto 0);
        ffc_macro_rst   : in     vl_logic;
        ffc_macropdb    : in     vl_logic;
        ffc_pcie_det_en : in     vl_logic_vector(1 downto 0);
        ffc_pcie_ct     : in     vl_logic_vector(1 downto 0);
        ffc_pfifo_clr   : in     vl_logic_vector(1 downto 0);
        ffc_dual_rst    : in     vl_logic;
        ffc_rrst        : in     vl_logic_vector(1 downto 0);
        ffc_rxpwdnb     : in     vl_logic_vector(1 downto 0);
        ffc_sb_inv_rx   : in     vl_logic_vector(1 downto 0);
        ffc_sb_pfifo_lp : in     vl_logic_vector(1 downto 0);
        ffc_signal_detect: in     vl_logic_vector(1 downto 0);
        ffc_sync_toggle : in     vl_logic;
        ffc_trst        : in     vl_logic;
        ffc_txpwdnb     : in     vl_logic_vector(1 downto 0);
        ffc_rx_div11_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_div11_mode: in     vl_logic_vector(1 downto 0);
        ffc_rx_rate_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_rate_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_gear_mode: in     vl_logic_vector(1 downto 0);
        ffc_rx_gear_mode: in     vl_logic_vector(1 downto 0);
        ffc_ldr_core2tx_en: in     vl_logic_vector(1 downto 0);
        ldr_core2tx     : in     vl_logic_vector(1 downto 0);
        ldr_core2tx_sd  : out    vl_logic_vector(1 downto 0);
        mc1_chif_ctl_ch0: in     vl_logic_vector(263 downto 0);
        mc1_chif_ctl_ch1: in     vl_logic_vector(263 downto 0);
        mc1_dif_ctl     : in     vl_logic_vector(159 downto 0);
        mc1_ser_ctl_ch0 : in     vl_logic_vector(87 downto 0);
        mc1_ser_ctl_ch1 : in     vl_logic_vector(87 downto 0);
        mc1_ser_ctl_dl  : in     vl_logic_vector(71 downto 0);
        pci_connect     : in     vl_logic_vector(1 downto 0);
        ffs_pcie_done   : out    vl_logic_vector(1 downto 0);
        ffs_pcie_con    : out    vl_logic_vector(1 downto 0);
        ff_tx_pclk      : out    vl_logic_vector(1 downto 0);
        ff_rx_pclk      : out    vl_logic_vector(1 downto 0);
        refck2core      : out    vl_logic;
        ffc_ck_core_rx  : in     vl_logic_vector(1 downto 0);
        ffc_ck_core_tx  : in     vl_logic;
        refc2core       : in     vl_logic;
        ck_core_rx      : out    vl_logic_vector(1 downto 0);
        ck_core_tx      : out    vl_logic;
        tck_aux_full    : in     vl_logic;
        plol            : in     vl_logic;
        rlol            : in     vl_logic_vector(1 downto 0);
        rlos            : in     vl_logic_vector(1 downto 0);
        pci_det_done    : in     vl_logic_vector(1 downto 0);
        reg2fpga_out_sd : in     vl_logic;
        ffs_plol        : out    vl_logic;
        ffs_rlol        : out    vl_logic_vector(1 downto 0);
        ffs_rlos        : out    vl_logic_vector(1 downto 0);
        reg2fpga_out    : out    vl_logic;
        rx_d_sd_0       : in     vl_logic_vector(9 downto 0);
        rx_d_sd_1       : in     vl_logic_vector(9 downto 0);
        sciaddr         : in     vl_logic_vector(5 downto 0);
        scienaux        : in     vl_logic;
        sciench0        : in     vl_logic;
        sciench1        : in     vl_logic;
        scird           : in     vl_logic;
        sciselaux       : in     vl_logic;
        sciselch0       : in     vl_logic;
        sciselch1       : in     vl_logic;
        sciwdata        : in     vl_logic_vector(7 downto 0);
        sciwstn         : in     vl_logic;
        rxr_clk_sd      : in     vl_logic_vector(1 downto 0);
        txp_clk_sd      : in     vl_logic_vector(1 downto 0);
        ser_sts_1_dl_25 : in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_0: in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27_1: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_0: in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28_1: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_0: in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29_1: in     vl_logic_vector(7 downto 0);
        ib_pwdnb        : out    vl_logic;
        txpll_pwdnb     : out    vl_logic;
        refck_pwdnb     : out    vl_logic;
        disable_dcu     : in     vl_logic;
        done_cfg        : in     vl_logic;
        scan_in         : in     vl_logic_vector(7 downto 0);
        scan_enable     : in     vl_logic;
        scan_reset      : in     vl_logic;
        scan_mode       : in     vl_logic;
        cout            : out    vl_logic_vector(19 downto 0);
        ff_rx_d_0       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_1       : out    vl_logic_vector(23 downto 0);
        ff_rx_f_clk     : out    vl_logic_vector(1 downto 0);
        ff_rx_h_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_f_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_h_clk     : out    vl_logic_vector(1 downto 0);
        pci_det_en      : out    vl_logic_vector(1 downto 0);
        ffs_cc_overrun  : out    vl_logic_vector(1 downto 0);
        ffs_cc_underrun : out    vl_logic_vector(1 downto 0);
        ffs_ls_sync_status: out    vl_logic_vector(1 downto 0);
        ffs_rxfbfifo_error: out    vl_logic_vector(1 downto 0);
        ffs_txfbfifo_error: out    vl_logic_vector(1 downto 0);
        ffs_skp_added   : out    vl_logic_vector(1 downto 0);
        ffs_skp_deleted : out    vl_logic_vector(1 downto 0);
        macrorst        : out    vl_logic;
        macropdb        : out    vl_logic;
        pcie_mode       : out    vl_logic_vector(1 downto 0);
        tx_d_sd_0       : out    vl_logic_vector(9 downto 0);
        tx_d_sd_1       : out    vl_logic_vector(9 downto 0);
        sciint          : out    vl_logic;
        scirdata        : out    vl_logic_vector(7 downto 0);
        ser_ctl_1_dl_0a : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_dl_0b : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_dl_0c : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_dl_0d : out    vl_logic_vector(7 downto 0);
        ser_ctl_5_dl_0e : out    vl_logic_vector(7 downto 0);
        ser_ctl_6_dl_12 : out    vl_logic_vector(7 downto 0);
        ser_ctl_7_dl_13 : out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_1_ch_10_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_8_ch_17_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_8_ch_17_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_9_ch_18_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_9_ch_18_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_10_ch_19_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_10_ch_19_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_11_ch_1a_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_11_ch_1a_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_12_ch_1b_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_12_ch_1b_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_13_ch_1c_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_13_ch_1c_1: out    vl_logic_vector(7 downto 0);
        ser_ctl_14_ch_1d_0: out    vl_logic_vector(7 downto 0);
        ser_ctl_14_ch_1d_1: out    vl_logic_vector(7 downto 0);
        sync_pulse      : out    vl_logic;
        rrst            : out    vl_logic_vector(1 downto 0);
        trst            : out    vl_logic;
        pci_det_ct      : out    vl_logic_vector(1 downto 0);
        pci_ei_en       : out    vl_logic_vector(1 downto 0);
        cdr_en_bitslip  : out    vl_logic_vector(1 downto 0);
        cfg_clk         : in     vl_logic;
        txpll_lol_from_nd: in     vl_logic;
        txpll_lol_to_nd : out    vl_logic;
        ffc_cdr_en_bitslip: in     vl_logic_vector(1 downto 0);
        ldr_rx2core_sd  : in     vl_logic_vector(1 downto 0);
        ldr_rx2core     : out    vl_logic_vector(1 downto 0);
        ser_mem_ch0     : out    vl_logic_vector(87 downto 0);
        ser_mem_ch1     : out    vl_logic_vector(87 downto 0);
        ser_mem_dl      : out    vl_logic_vector(71 downto 0);
        scan_out        : out    vl_logic_vector(7 downto 0);
        bs2pad          : out    vl_logic_vector(1 downto 0);
        bs4pad          : in     vl_logic_vector(1 downto 0);
        bs4refclk       : in     vl_logic;
        shift_dr        : in     vl_logic;
        si_jtag         : in     vl_logic;
        clock_dr_in     : in     vl_logic;
        update_dr       : in     vl_logic;
        mode_jtag       : in     vl_logic_vector(1 downto 0);
        rst_jtag        : in     vl_logic;
        so_jtag         : out    vl_logic;
        clock_dr_out    : out    vl_logic;
        shiftdrn_out    : out    vl_logic;
        updatedr_out    : out    vl_logic;
        mode_jtag_sd    : out    vl_logic
    );
end pcs_dual;
