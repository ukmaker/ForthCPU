library verilog;
use verilog.vl_types.all;
entity vhiv1s is
    port(
        Z               : out    vl_logic
    );
end vhiv1s;
