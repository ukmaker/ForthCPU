library verilog;
use verilog.vl_types.all;
entity sbnx2v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end sbnx2v1s;
