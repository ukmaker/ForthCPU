library verilog;
use verilog.vl_types.all;
entity delc12 is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end delc12;
