library verilog;
use verilog.vl_types.all;
entity pcs_aoi22_2 is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        X               : out    vl_logic
    );
end pcs_aoi22_2;
