library verilog;
use verilog.vl_types.all;
entity dcu_top is
    port(
        hdinn0          : in     vl_logic;
        hdinn1          : in     vl_logic;
        hdinp0          : in     vl_logic;
        hdinp1          : in     vl_logic;
        iref_50urpoly   : in     vl_logic_vector(1 downto 0);
        iref_50uconst   : in     vl_logic_vector(1 downto 0);
        ffc_cdr_en_bitslip: in     vl_logic_vector(1 downto 0);
        ffc_ck_core_rx  : in     vl_logic_vector(1 downto 0);
        ffc_ck_core_tx  : in     vl_logic;
        txbit_clkp_from_nd: in     vl_logic;
        txbit_clkn_from_nd: in     vl_logic;
        refck_from_ndp  : in     vl_logic;
        refck_from_ndn  : in     vl_logic;
        refclkn         : in     vl_logic;
        refclkp         : in     vl_logic;
        sync_ndp        : in     vl_logic;
        sync_ndn        : in     vl_logic;
        cin             : in     vl_logic_vector(11 downto 0);
        ff_ebrd_clk     : in     vl_logic_vector(1 downto 0);
        ff_rxi_clk      : in     vl_logic_vector(1 downto 0);
        ff_tx_d_0       : in     vl_logic_vector(23 downto 0);
        ff_tx_d_1       : in     vl_logic_vector(23 downto 0);
        ff_txi_clk      : in     vl_logic_vector(1 downto 0);
        ffc_ei_en       : in     vl_logic_vector(1 downto 0);
        ffc_enable_cgalign: in     vl_logic_vector(1 downto 0);
        ffc_fb_loopback : in     vl_logic_vector(1 downto 0);
        ffc_tx_lane_rst : in     vl_logic_vector(1 downto 0);
        ffc_rx_lane_rst : in     vl_logic_vector(1 downto 0);
        ffc_macro_rst   : in     vl_logic;
        ffc_pcie_det_en : in     vl_logic_vector(1 downto 0);
        ffc_pcie_ct     : in     vl_logic_vector(1 downto 0);
        ffc_pfifo_clr   : in     vl_logic_vector(1 downto 0);
        ffc_macropdb    : in     vl_logic;
        ffc_dual_rst    : in     vl_logic;
        ffc_rrst        : in     vl_logic_vector(1 downto 0);
        ffc_rpwdnb      : in     vl_logic_vector(1 downto 0);
        ffc_sb_inv_rx   : in     vl_logic_vector(1 downto 0);
        ffc_sb_pfifo_lp : in     vl_logic_vector(1 downto 0);
        ffc_signal_detect: in     vl_logic_vector(1 downto 0);
        ffc_sync_toggle : in     vl_logic;
        ffc_trst        : in     vl_logic;
        ffc_tpwdnb      : in     vl_logic_vector(1 downto 0);
        ffc_rx_div11_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_div11_mode: in     vl_logic_vector(1 downto 0);
        ffc_rx_rate_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_rate_mode: in     vl_logic_vector(1 downto 0);
        ffc_tx_gear_mode: in     vl_logic_vector(1 downto 0);
        ffc_rx_gear_mode: in     vl_logic_vector(1 downto 0);
        ffc_ldr_core2tx_en: in     vl_logic_vector(1 downto 0);
        ldr_core2tx     : in     vl_logic_vector(1 downto 0);
        txpll_lol_from_nd: in     vl_logic;
        sciaddr         : in     vl_logic_vector(5 downto 0);
        scienaux        : in     vl_logic;
        sciench0        : in     vl_logic;
        sciench1        : in     vl_logic;
        scird           : in     vl_logic;
        sciselaux       : in     vl_logic;
        sciselch0       : in     vl_logic;
        sciselch1       : in     vl_logic;
        sciwdata        : in     vl_logic_vector(7 downto 0);
        sciwstn         : in     vl_logic;
        cyawstn         : in     vl_logic;
        cfg_clk         : in     vl_logic;
        done_cfg        : in     vl_logic;
        shift_dr        : in     vl_logic;
        si_jtag         : in     vl_logic;
        clock_dr_in     : in     vl_logic;
        update_dr       : in     vl_logic;
        mode_jtag       : in     vl_logic_vector(1 downto 0);
        rst_jtag        : in     vl_logic;
        scan_in         : in     vl_logic_vector(7 downto 0);
        scan_enable     : in     vl_logic;
        scan_reset      : in     vl_logic;
        scan_mode       : in     vl_logic;
        mc1_chif_ctl_ch0: in     vl_logic_vector(263 downto 0);
        mc1_chif_ctl_ch1: in     vl_logic_vector(263 downto 0);
        mc1_dif_ctl     : in     vl_logic_vector(159 downto 0);
        mc1_ser_ctl_ch0 : in     vl_logic_vector(87 downto 0);
        mc1_ser_ctl_ch1 : in     vl_logic_vector(87 downto 0);
        mc1_ser_ctl_dl  : in     vl_logic_vector(71 downto 0);
        disable_dcu     : in     vl_logic;
        txbit_clkp_to_nd: out    vl_logic;
        txbit_clkn_to_nd: out    vl_logic;
        hdoutn0         : out    vl_logic;
        hdoutn1         : out    vl_logic;
        hdoutp0         : out    vl_logic;
        hdoutp1         : out    vl_logic;
        atstp           : inout  vl_logic;
        atstn           : inout  vl_logic;
        ffs_pcie_con    : out    vl_logic_vector(1 downto 0);
        ffs_pcie_done   : out    vl_logic_vector(1 downto 0);
        ffs_plol        : out    vl_logic;
        ffs_rlol        : out    vl_logic_vector(1 downto 0);
        ffs_rlos        : out    vl_logic_vector(1 downto 0);
        refck2core      : out    vl_logic;
        ff_rx_pclk      : out    vl_logic_vector(1 downto 0);
        ff_tx_pclk      : out    vl_logic_vector(1 downto 0);
        refck2ndp       : out    vl_logic;
        refck2ndn       : out    vl_logic;
        reg2fpga_out    : out    vl_logic;
        sync2ndp        : out    vl_logic;
        sync2ndn        : out    vl_logic;
        cout            : out    vl_logic_vector(19 downto 0);
        ff_rx_d_0       : out    vl_logic_vector(23 downto 0);
        ff_rx_d_1       : out    vl_logic_vector(23 downto 0);
        ff_rx_f_clk     : out    vl_logic_vector(1 downto 0);
        ff_rx_h_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_f_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_h_clk     : out    vl_logic_vector(1 downto 0);
        ffs_cc_overrun  : out    vl_logic_vector(1 downto 0);
        ffs_cc_underrun : out    vl_logic_vector(1 downto 0);
        ffs_ls_sync_status: out    vl_logic_vector(1 downto 0);
        ffs_rxfbfifo_error: out    vl_logic_vector(1 downto 0);
        ffs_txfbfifo_error: out    vl_logic_vector(1 downto 0);
        ffs_skp_added   : out    vl_logic_vector(1 downto 0);
        ffs_skp_deleted : out    vl_logic_vector(1 downto 0);
        ldr_rx2core     : out    vl_logic_vector(1 downto 0);
        txpll_lol_to_nd : out    vl_logic;
        sciint          : out    vl_logic;
        scirdata        : out    vl_logic_vector(7 downto 0);
        so_jtag         : out    vl_logic;
        clock_dr_out    : out    vl_logic;
        shiftdrn_out    : out    vl_logic;
        updatedr_out    : out    vl_logic;
        scan_out        : out    vl_logic_vector(7 downto 0);
        vcca            : inout  vl_logic;
        vcca25          : inout  vl_logic;
        vccatx0         : inout  vl_logic;
        vccatx1         : inout  vl_logic;
        vccarx0         : inout  vl_logic;
        vccarx1         : inout  vl_logic;
        vcchtx0         : inout  vl_logic;
        vcchtx1         : inout  vl_logic;
        vcchrx0         : inout  vl_logic;
        vcchrx1         : inout  vl_logic;
        vssa            : inout  vl_logic;
        vssach0         : inout  vl_logic;
        vssach1         : inout  vl_logic
    );
end dcu_top;
