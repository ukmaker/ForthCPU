library verilog;
use verilog.vl_types.all;
entity pcs_channel_top is
    port(
        bus8bit_sel     : in     vl_logic;
        bist_rx_data_sel: in     vl_logic;
        char_test_data  : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic;
        ebrd_clk        : in     vl_logic;
        fbw_clk         : in     vl_logic;
        ff_tx_d         : in     vl_logic_vector(23 downto 0);
        ffc_ei_en       : in     vl_logic;
        ffc_enable_cgalign: in     vl_logic;
        ffc_fb_loopback : in     vl_logic;
        ffc_pcie_det_en : in     vl_logic;
        ffc_pcie_ct     : in     vl_logic;
        pfifor_clr      : in     vl_logic;
        pfifow_clr      : in     vl_logic;
        pfifo_clr_sel   : in     vl_logic;
        ffc_rxpwdnb     : in     vl_logic;
        ffc_rx_div11_mode: in     vl_logic;
        ffc_tx_div11_mode: in     vl_logic;
        ffc_rx_rate_mode: in     vl_logic;
        ffc_tx_rate_mode: in     vl_logic;
        ffc_rx_gear_mode: in     vl_logic;
        ffc_tx_gear_mode: in     vl_logic;
        ffc_cdr_en_bitslip: in     vl_logic;
        ffc_sb_inv_rx   : in     vl_logic;
        ffc_sb_pfifo_lp : in     vl_logic;
        ffc_signal_detect: in     vl_logic;
        ffc_txpwdnb     : in     vl_logic;
        rxf_clk         : in     vl_logic;
        txf_clk         : in     vl_logic;
        fmbist_data     : in     vl_logic_vector(9 downto 0);
        force_int       : in     vl_logic;
        ffc_ldr_core2tx_en: in     vl_logic;
        mc1_chif_ctl    : in     vl_logic_vector(263 downto 0);
        mc1_ser_ctl     : in     vl_logic_vector(87 downto 0);
        pci_connect     : in     vl_logic;
        pcie_rxpolarity : in     vl_logic;
        pcie_txcompliance: in     vl_logic;
        pcie_txdetrx_pr2tlb: in     vl_logic;
        pcie_txelecidle : in     vl_logic;
        pcs_ctl_3_dl_02 : in     vl_logic_vector(7 downto 0);
        plol            : in     vl_logic;
        rstb_txf        : in     vl_logic;
        rstb_txp        : in     vl_logic;
        rstb_ebrd       : in     vl_logic;
        rstb_rxr        : in     vl_logic;
        rstb_fbw        : in     vl_logic;
        rstb_rxf        : in     vl_logic;
        rxr_clk         : in     vl_logic;
        done_cfg        : in     vl_logic;
        reg_load        : in     vl_logic;
        goe_r2          : in     vl_logic;
        goe_load        : in     vl_logic;
        sciaddr         : in     vl_logic_vector(5 downto 0);
        sciwdata        : in     vl_logic_vector(7 downto 0);
        scird           : in     vl_logic;
        cyawstn         : in     vl_logic;
        sciench         : in     vl_logic;
        sciselch        : in     vl_logic;
        ser_sts_1_ch_26 : in     vl_logic_vector(7 downto 0);
        ser_sts_2_ch_27 : in     vl_logic_vector(7 downto 0);
        ser_sts_3_ch_28 : in     vl_logic_vector(7 downto 0);
        ser_sts_4_ch_29 : in     vl_logic_vector(7 downto 0);
        serdes_rxd      : in     vl_logic_vector(9 downto 0);
        txp_clk         : in     vl_logic;
        xge_mode        : in     vl_logic;
        ff_rx_d         : out    vl_logic_vector(23 downto 0);
        pci_det_en      : out    vl_logic;
        ffs_cc_overrun  : out    vl_logic;
        ffs_cc_underrun : out    vl_logic;
        ffs_ls_sync_status: out    vl_logic;
        ffs_rxfbfifo_error: out    vl_logic;
        ffs_txfbfifo_error: out    vl_logic;
        pcie_mode       : out    vl_logic;
        pcie_phystatus  : out    vl_logic;
        pcie_rxvalid    : out    vl_logic;
        skp_add         : out    vl_logic;
        skp_del         : out    vl_logic;
        pfifo_error     : out    vl_logic;
        full_d          : out    vl_logic;
        empty_d         : out    vl_logic;
        scirdata_01     : out    vl_logic_vector(7 downto 0);
        sciint_10       : out    vl_logic;
        rx_ch           : out    vl_logic;
        txd_sd          : out    vl_logic_vector(9 downto 0);
        ser_ctl_1_ch_10 : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_ch_11 : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_ch_12 : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_ch_13 : out    vl_logic_vector(7 downto 0);
        ser_ctl_5_ch_14 : out    vl_logic_vector(7 downto 0);
        ser_ctl_6_ch_15 : out    vl_logic_vector(7 downto 0);
        ser_ctl_7_ch_16 : out    vl_logic_vector(7 downto 0);
        ser_ctl_8_ch_17 : out    vl_logic_vector(7 downto 0);
        ser_ctl_9_ch_18 : out    vl_logic_vector(7 downto 0);
        ser_ctl_10_ch_19: out    vl_logic_vector(7 downto 0);
        ser_ctl_11_ch_1a: out    vl_logic_vector(7 downto 0);
        ser_ctl_12_ch_1b: out    vl_logic_vector(7 downto 0);
        ser_ctl_13_ch_1c: out    vl_logic_vector(7 downto 0);
        ser_ctl_14_ch_1d: out    vl_logic_vector(7 downto 0);
        rst_ctl_1_ch_1f : out    vl_logic_vector(7 downto 0);
        pcs_ctl_3_ch_02 : out    vl_logic_vector(7 downto 0);
        tobist_data     : out    vl_logic_vector(9 downto 0);
        pci_det_ct      : out    vl_logic;
        pci_ei_en       : out    vl_logic;
        cdr_en_bitslip  : out    vl_logic;
        ser_mem         : out    vl_logic_vector(87 downto 0)
    );
end pcs_channel_top;
