library verilog;
use verilog.vl_types.all;
entity SEH_INV_S_6 is
    port(
        X               : out    vl_logic;
        A               : in     vl_logic
    );
end SEH_INV_S_6;
