library verilog;
use verilog.vl_types.all;
entity CDCHK_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end CDCHK_UDP;
