library verilog;
use verilog.vl_types.all;
entity NNP_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end NNP_UDP;
