library verilog;
use verilog.vl_types.all;
entity mem_top_reno is
    generic(
        CFG_ARRAY_ROW_COUNT: integer := 14;
        CFG_WORDWIDTH   : integer := 8;
        TRIM_ARRAY_ROW_COUNT: integer := 4;
        TRIM_WORDWIDTH  : integer := 8;
        FLUT_ARRAY_ROW_COUNT: integer := 16;
        FLUT_WORDWIDTH  : integer := 7;
        \CFG_SEL_ARRAY\ : integer := 16;
        \DONEBIT_SEL_ARRAY\: integer := 8;
        \FLUT_SEL_ARRAY\: integer := 4;
        I2CMSB_SEL_ARRAY: integer := 2;
        \TRIM_SEL_ARRAY\: integer := 1;
        CFG_EEPROM      : string  := "cfg_eeprom.hex";
        TRIM_EEPROM     : string  := "trim_eeprom.hex";
        FLUT_EEPROM     : string  := "flut_eeprom.hex";
        I2CADDRESS      : string  := "i2caddress.hex"
    );
    port(
        a_test_in       : in     vl_logic;
        a_test_out      : inout  vl_logic;
        a_vppout        : out    vl_logic;
        cfg_sel_array   : in     vl_logic;
        cfgtrim_drvmcbus: in     vl_logic;
        cfgtrim_load_addrlat: in     vl_logic;
        cfgtrim_load_datareg: in     vl_logic;
        cfgtrim_sel_datareg: in     vl_logic;
        data_enable     : in     vl_logic;
        donebit         : out    vl_logic;
        donebit_sel_array: in     vl_logic;
        d_test_out      : out    vl_logic;
        enable_erase    : in     vl_logic;
        enable_program  : in     vl_logic;
        faultlog_load_soft_datareg: in     vl_logic;
        faultlog_sel_twi: in     vl_logic;
        flut_col_addr   : in     vl_logic_vector(2 downto 0);
        flut_drvmcbus   : in     vl_logic;
        flut_load_datareg: in     vl_logic;
        flut_row_addr   : in     vl_logic_vector(3 downto 0);
        flut_sel_array  : in     vl_logic;
        flut_sel_sdatareg: in     vl_logic;
        hvblock         : in     vl_logic;
        i2csa           : out    vl_logic_vector(6 downto 3);
        i2csa_done      : out    vl_logic;
        i2csa_drvmcbus  : in     vl_logic;
        i2csa_load_datareg: in     vl_logic;
        i2csa_lsb       : in     vl_logic_vector(2 downto 0);
        i2csa_sel_array : in     vl_logic;
        iabias_25u      : inout  vl_logic;
        ibgtrim_reg     : in     vl_logic_vector(2 downto 0);
        ihvout0_n5u     : inout  vl_logic;
        ihvout1_n5u     : inout  vl_logic;
        ihvout2_n5u     : inout  vl_logic;
        ihvout3_n5u     : inout  vl_logic;
        ii2c_25u        : inout  vl_logic;
        ioa_25u         : inout  vl_logic;
        iosc_25u        : inout  vl_logic;
        irefpad_bot_n10u: inout  vl_logic;
        irefpad_top_n10u: inout  vl_logic;
        mcbus_data      : inout  vl_logic_vector(7 downto 0);
        mfg_cfgsel      : in     vl_logic;
        mfg_dbg_iref    : in     vl_logic;
        mfg_dbg_vref    : in     vl_logic;
        mfg_donesel     : in     vl_logic;
        mfg_faultsel    : in     vl_logic;
        mfg_i2csel      : in     vl_logic;
        mfg_mcgforce    : in     vl_logic;
        mfg_mcgoe       : in     vl_logic;
        mfg_progallrows : in     vl_logic;
        mfg_progoddeve  : in     vl_logic;
        mfg_trimsel     : in     vl_logic;
        mfg_vhien       : in     vl_logic;
        mfg_vppdiv      : in     vl_logic;
        mfg_vppen       : in     vl_logic;
        mfg_vppoe       : in     vl_logic;
        mfg_vpp_pf      : in     vl_logic;
        por_n           : in     vl_logic;
        slrtrim_reg     : in     vl_logic_vector(2 downto 0);
        trim_sel_array  : in     vl_logic;
        twi_data        : in     vl_logic_vector(7 downto 0);
        v2p1            : in     vl_logic;
        vbgtrim_reg     : in     vl_logic_vector(2 downto 0);
        vdbg            : inout  vl_logic;
        vddd            : in     vl_logic;
        vhi             : out    vl_logic;
        vppoff          : out    vl_logic;
        vpptrim_erase   : in     vl_logic_vector(4 downto 0);
        vpptrim_program : in     vl_logic_vector(4 downto 0);
        vssd            : in     vl_logic
    );
end mem_top_reno;
