library verilog;
use verilog.vl_types.all;
entity jtag_logic is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 1;
        DECRYPTION      : integer := 1
    );
    port(
        jsel_byp        : out    vl_logic;
        jsel_cfg        : out    vl_logic;
        jsel_sec        : out    vl_logic;
        jsel_com        : out    vl_logic;
        jsel_com_lsbf   : out    vl_logic;
        jsel_com_msbf   : out    vl_logic;
        jcap_com_word4  : out    vl_logic;
        jshf_com_byte1  : out    vl_logic;
        jshf_com_byte1_msbf: out    vl_logic;
        jshf_com_byte2  : out    vl_logic;
        jshf_com_byte4  : out    vl_logic;
        jshf_com_byte8  : out    vl_logic;
        jshf_com_byte9_msbf: out    vl_logic;
        jshf_com_word4  : out    vl_logic;
        jshf_com_word4_msbf: out    vl_logic;
        jbuf8_s01       : out    vl_logic;
        jbuf8_p08       : out    vl_logic;
        jbuf8_rst       : out    vl_logic;
        jsel_busy       : out    vl_logic;
        jsel_er1        : out    vl_logic;
        jsel_er2        : out    vl_logic;
        jsel_bsr        : out    vl_logic;
        jsel_sram_asr   : out    vl_logic;
        jsel_dsr        : out    vl_logic;
        jsel_mfg        : out    vl_logic;
        jsel_iscan      : out    vl_logic;
        jsel_extspi_i   : out    vl_logic;
        jsel_extspi     : out    vl_logic;
        lsc_iscan_m     : out    vl_logic_vector(7 downto 0);
        iscan_en        : out    vl_logic_vector(7 downto 0);
        test_mode_i     : out    vl_logic;
        non_test_mode_i : out    vl_logic;
        j_enable_qual   : out    vl_logic;
        j_enable_x_qual : out    vl_logic;
        j_disable_qual  : out    vl_logic;
        rti2d           : out    vl_logic;
        bsrclk          : out    vl_logic;
        shiftdr_bs      : out    vl_logic;
        updatedr_bs     : out    vl_logic;
        bsmode1         : out    vl_logic;
        bsmode2         : out    vl_logic;
        bsmode3         : out    vl_logic;
        ac_mode         : out    vl_logic;
        ac_test         : out    vl_logic;
        ac_clear        : out    vl_logic;
        tsall_ctrl      : out    vl_logic;
        isptcy_rtier1   : out    vl_logic;
        isptcy_rtier2   : out    vl_logic;
        isptcy_shcap    : out    vl_logic;
        isptcy_update   : out    vl_logic;
        isptcy_ener1    : out    vl_logic;
        isptcy_ener2    : out    vl_logic;
        isptcy_resetb   : out    vl_logic;
        isptcy_tdi      : out    vl_logic;
        lsc_read_status_m: out    vl_logic;
        lsc_read_mfg_status_m: out    vl_logic;
        lsc_read_pes_m  : out    vl_logic;
        lsc_read_mes_m  : out    vl_logic;
        lsc_read_hes_m  : out    vl_logic;
        lsc_read_trim_m : out    vl_logic;
        lsc_read_comp_dic_m: out    vl_logic;
        lsc_prog_pes_m  : out    vl_logic;
        lsc_prog_mes_m  : out    vl_logic;
        lsc_prog_hes_m  : out    vl_logic;
        lsc_prog_trim_m : out    vl_logic;
        jexit_fl_offline: out    vl_logic;
        jexit_normal    : out    vl_logic;
        jtag_active     : out    vl_logic;
        tdrclk_sw_i     : out    vl_logic;
        jenable_tran    : out    vl_logic;
        jenable_offl    : out    vl_logic;
        jrst_isc_done_i : out    vl_logic;
        jset_isc_done_i : out    vl_logic;
        jaccess_sram    : out    vl_logic;
        jaccess_flash   : out    vl_logic;
        jaccess_fl_norm : out    vl_logic;
        jaccess_fl_sudo : out    vl_logic;
        jaccess_fl_safe : out    vl_logic;
        jaccess_efuse   : out    vl_logic;
        jaccess_ef_norm : out    vl_logic;
        jaccess_ef_sudo : out    vl_logic;
        jaccess_ef_safe : out    vl_logic;
        jaccess_tag     : out    vl_logic;
        jaccess_flash_all: out    vl_logic;
        ins_dsr_1bit    : out    vl_logic;
        ins_dsr_1byte   : out    vl_logic;
        jburst_pause    : out    vl_logic;
        jburst_01       : out    vl_logic;
        jburst_08       : out    vl_logic;
        j_ins_prog_com  : out    vl_logic;
        jburst_en       : out    vl_logic;
        jpspi_en_norm   : out    vl_logic;
        jpspi_en_stack  : out    vl_logic;
        jpspi_en_int    : out    vl_logic;
        jpspi_param     : out    vl_logic_vector(7 downto 0);
        por             : in     vl_logic;
        tck             : in     vl_logic;
        tms             : in     vl_logic;
        tdi             : in     vl_logic;
        tlreset         : in     vl_logic;
        rti_r           : in     vl_logic;
        seldr_ss        : in     vl_logic;
        capdr_ss        : in     vl_logic;
        shiftdr_ss      : in     vl_logic;
        updr_ss         : in     vl_logic;
        exit1dr_ss      : in     vl_logic;
        exit2dr_ss      : in     vl_logic;
        ShiftDR         : in     vl_logic;
        UpdateDR        : in     vl_logic;
        ClockDR         : in     vl_logic;
        jconfig_dat     : in     vl_logic_vector(3 downto 0);
        mfg_prog_sel    : in     vl_logic_vector(3 downto 0);
        mfg_iscan_sel   : in     vl_logic_vector(2 downto 0);
        mfg_iscan_en    : in     vl_logic;
        mfg_pshf_sel    : in     vl_logic;
        jpspi_ctrl      : in     vl_logic_vector(15 downto 0);
        extest_i        : in     vl_logic;
        extest_pulse_i  : in     vl_logic;
        extest_train_i  : in     vl_logic;
        intest_i        : in     vl_logic;
        clamp_i         : in     vl_logic;
        highz_i         : in     vl_logic;
        sample_prld_i   : in     vl_logic;
        bypass_i        : in     vl_logic;
        verify_id_i     : in     vl_logic;
        idcode_pub_i    : in     vl_logic;
        uidcode_pub_i   : in     vl_logic;
        usercode_i      : in     vl_logic;
        read_temp_i     : in     vl_logic;
        lsc_device_ctrl_i: in     vl_logic;
        lsc_shift_password_i: in     vl_logic;
        lsc_read_status_i: in     vl_logic;
        lsc_check_busy_i: in     vl_logic;
        lsc_refresh_i   : in     vl_logic;
        lsc_bitstream_burst_i: in     vl_logic;
        lsc_i2ci_crbr_wt_i: in     vl_logic;
        lsc_i2ci_txdr_wt_i: in     vl_logic;
        lsc_i2ci_rxdr_rd_i: in     vl_logic;
        lsc_i2ci_sr_rd_i: in     vl_logic;
        ip_a_i          : in     vl_logic;
        ip_b_i          : in     vl_logic;
        iptest_a_i      : in     vl_logic;
        iptest_b_i      : in     vl_logic;
        lsc_prog_spi_i  : in     vl_logic;
        idcode_prv_i    : in     vl_logic;
        read_pes_i      : in     vl_logic;
        mfg_shift_i     : in     vl_logic;
        isc_enable_i    : in     vl_logic;
        isc_enable_x_i  : in     vl_logic;
        isc_disable_i   : in     vl_logic;
        isc_program_i   : in     vl_logic;
        isc_noop_i      : in     vl_logic;
        isc_prog_ucode_i: in     vl_logic;
        isc_read_i      : in     vl_logic;
        isc_erase_i     : in     vl_logic;
        isc_discharge_i : in     vl_logic;
        isc_prog_done_i : in     vl_logic;
        isc_erase_done_i: in     vl_logic;
        isc_prog_sec_i  : in     vl_logic;
        isc_prog_secplus_i: in     vl_logic;
        isc_data_shift_i: in     vl_logic;
        isc_addr_shift_i: in     vl_logic;
        lsc_init_addr_i : in     vl_logic;
        lsc_write_addr_i: in     vl_logic;
        lsc_prog_incr_rti_i: in     vl_logic;
        lsc_prog_incr_enc_i: in     vl_logic;
        lsc_prog_incr_cmp_i: in     vl_logic;
        lsc_prog_incr_cne_i: in     vl_logic;
        lsc_vfy_incr_rti_i: in     vl_logic;
        lsc_prog_ctrl0_i: in     vl_logic;
        lsc_read_ctrl0_i: in     vl_logic;
        lsc_reset_crc_i : in     vl_logic;
        lsc_read_crc_i  : in     vl_logic;
        lsc_prog_sed_crc_i: in     vl_logic;
        lsc_read_sed_crc_i: in     vl_logic;
        lsc_prog_password_i: in     vl_logic;
        lsc_read_password_i: in     vl_logic;
        lsc_prog_cipher_key_i: in     vl_logic;
        lsc_read_cipher_key_i: in     vl_logic;
        lsc_prog_feature_i: in     vl_logic;
        lsc_read_feature_i: in     vl_logic;
        lsc_prog_feabits_i: in     vl_logic;
        lsc_read_feabits_i: in     vl_logic;
        lsc_prog_otps_i : in     vl_logic;
        lsc_read_otps_i : in     vl_logic;
        lsc_write_comp_dic_i: in     vl_logic;
        lsc_write_bus_addr_i: in     vl_logic;
        lsc_pcs_write_i : in     vl_logic;
        lsc_pcs_read_i  : in     vl_logic;
        lsc_ebr_write_i : in     vl_logic;
        lsc_ebr_read_i  : in     vl_logic;
        lsc_prog_incr_nv_i: in     vl_logic;
        lsc_read_incr_nv_i: in     vl_logic;
        lsc_init_addr_ufm_i: in     vl_logic;
        lsc_prog_tag_i  : in     vl_logic;
        lsc_erase_tag_i : in     vl_logic;
        lsc_read_tag_i  : in     vl_logic;
        lsc_prog_pes_i  : in     vl_logic;
        lsc_mtest_i     : in     vl_logic;
        lsc_mtrim_i     : in     vl_logic;
        lsc_mdata_i     : in     vl_logic;
        lsc_iscan_i     : in     vl_logic;
        mfg_en          : in     vl_logic;
        mc1_er1_exist   : in     vl_logic;
        mc1_er2_exist   : in     vl_logic;
        isc_enabled     : in     vl_logic;
        isc_done        : in     vl_logic;
        isc_disable_completing: in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic
    );
end jtag_logic;
