library verilog;
use verilog.vl_types.all;
entity SEH_AOI22_S_4 is
    port(
        X               : out    vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic
    );
end SEH_AOI22_S_4;
