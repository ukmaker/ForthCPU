library verilog;
use verilog.vl_types.all;
entity ser_rx_misc is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end ser_rx_misc;
