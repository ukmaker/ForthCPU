library verilog;
use verilog.vl_types.all;
entity njtag_logic is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 1;
        DECRYPTION      : integer := 1
    );
    port(
        njsel_byp       : out    vl_logic;
        njsel_cfg       : out    vl_logic;
        njsel_sec       : out    vl_logic;
        njsel_dsr       : out    vl_logic;
        njsel_com       : out    vl_logic;
        njcap_com_word4_norm: out    vl_logic;
        njcap_com_word4_slow: out    vl_logic;
        njshf_com_byte1 : out    vl_logic;
        njshf_com_byte2 : out    vl_logic;
        njshf_com_byte4 : out    vl_logic;
        njshf_com_byte8 : out    vl_logic;
        njshf_com_byte9 : out    vl_logic;
        njshf_com_word4 : out    vl_logic;
        njsel_extspi    : out    vl_logic;
        nj_cmd_read_dat : out    vl_logic;
        nj_enable_qual  : out    vl_logic;
        nj_enable_x_qual: out    vl_logic;
        nj_disable_qual : out    vl_logic;
        bse_end_cqual   : out    vl_logic;
        nj_check_crc    : out    vl_logic;
        nj_exec_a       : out    vl_logic;
        nj_exec_b       : out    vl_logic;
        nj_exec_c       : out    vl_logic;
        nj_exec_d       : out    vl_logic;
        nj_exec_e       : out    vl_logic;
        nj_exec_f       : out    vl_logic;
        njexit_fl_offline: out    vl_logic;
        njexit_normal   : out    vl_logic;
        njtag_active    : out    vl_logic;
        njtag_active_nsed: out    vl_logic;
        njenable_tran   : out    vl_logic;
        njenable_offl   : out    vl_logic;
        njrst_isc_done_c: out    vl_logic;
        njset_isc_done_c: out    vl_logic;
        njaccess_sram   : out    vl_logic;
        njaccess_flash  : out    vl_logic;
        njaccess_fl_norm: out    vl_logic;
        njaccess_fl_sudo: out    vl_logic;
        njaccess_fl_safe: out    vl_logic;
        njaccess_efuse  : out    vl_logic;
        njaccess_ef_norm: out    vl_logic;
        njaccess_ef_sudo: out    vl_logic;
        njaccess_ef_safe: out    vl_logic;
        njaccess_tag    : out    vl_logic;
        njaccess_flash_all: out    vl_logic;
        njtag_bse_en    : out    vl_logic;
        njtag_slv_en    : out    vl_logic;
        nj_cmd_ndata    : out    vl_logic;
        nj_cmd_read     : out    vl_logic;
        nj_cmd_incr     : out    vl_logic;
        nj_cmd_prog     : out    vl_logic;
        nj_cmd_prog_incr: out    vl_logic;
        nj_cmd_read_incr: out    vl_logic;
        nj_cmd_prog_dsr : out    vl_logic;
        nj_cmd_read_dsr : out    vl_logic;
        nj_cmd_read_com : out    vl_logic;
        nj_cmd_prog_com : out    vl_logic;
        nj_cmd_read_fslow: out    vl_logic;
        sed_cmd_read_incr: out    vl_logic;
        njtag_data_byte : out    vl_logic_vector(15 downto 0);
        extra_dsr_cnt   : out    vl_logic;
        lsc_pcs_rw_c    : out    vl_logic;
        njm_invalid_c   : out    vl_logic;
        njr_invalid_c   : out    vl_logic;
        njs_invalid_c   : out    vl_logic;
        sed_invalid_c   : out    vl_logic;
        cmd_dsr_1byte   : out    vl_logic;
        njvfy_rst_exec  : out    vl_logic;
        njpspi_en_norm  : out    vl_logic;
        njpspi_en_stack : out    vl_logic;
        njpspi_en_int   : out    vl_logic;
        njpspi_param    : out    vl_logic_vector(7 downto 0);
        njburst_inp     : out    vl_logic;
        DSR_LENGTH      : in     vl_logic_vector(15 downto 0);
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        scanen          : in     vl_logic;
        jtag_active_smsync: in     vl_logic;
        p_scm           : in     vl_logic;
        njport_active   : in     vl_logic;
        njport_exec     : in     vl_logic;
        njshf_dum       : in     vl_logic;
        njbse_rxcmd     : in     vl_logic;
        njbse_rxdec     : in     vl_logic;
        sed_boot        : in     vl_logic;
        sed_en_adv      : in     vl_logic;
        njconfig_dat    : in     vl_logic_vector(3 downto 0);
        njshf_dat       : in     vl_logic;
        post_dec        : in     vl_logic;
        post_inf1       : in     vl_logic;
        post_inf2       : in     vl_logic;
        post_inf3       : in     vl_logic;
        post_crc        : in     vl_logic;
        fsm_exec_e      : in     vl_logic;
        fsm_exec_f      : in     vl_logic;
        njpspi_ctrl     : in     vl_logic_vector(15 downto 0);
        bypass_c        : in     vl_logic;
        verify_id_c     : in     vl_logic;
        idcode_pub_c    : in     vl_logic;
        uidcode_pub_c   : in     vl_logic;
        usercode_c      : in     vl_logic;
        read_temp_c     : in     vl_logic;
        lsc_device_ctrl_c: in     vl_logic;
        lsc_shift_password_c: in     vl_logic;
        lsc_read_status_c: in     vl_logic;
        lsc_check_busy_c: in     vl_logic;
        lsc_refresh_c   : in     vl_logic;
        lsc_bitstream_burst_c: in     vl_logic;
        lsc_i2ci_crbr_wt_c: in     vl_logic;
        lsc_i2ci_txdr_wt_c: in     vl_logic;
        lsc_i2ci_rxdr_rd_c: in     vl_logic;
        lsc_i2ci_sr_rd_c: in     vl_logic;
        lsc_prog_spi_c  : in     vl_logic;
        idcode_prv_c    : in     vl_logic;
        read_pes_c      : in     vl_logic;
        isc_enable_c    : in     vl_logic;
        isc_enable_x_c  : in     vl_logic;
        isc_disable_c   : in     vl_logic;
        isc_program_c   : in     vl_logic;
        isc_noop_c      : in     vl_logic;
        isc_prog_ucode_c: in     vl_logic;
        isc_read_c      : in     vl_logic;
        isc_erase_c     : in     vl_logic;
        isc_prog_done_c : in     vl_logic;
        isc_erase_done_c: in     vl_logic;
        isc_prog_sec_c  : in     vl_logic;
        isc_prog_secplus_c: in     vl_logic;
        isc_data_shift_c: in     vl_logic;
        isc_addr_shift_c: in     vl_logic;
        lsc_init_addr_c : in     vl_logic;
        lsc_write_addr_c: in     vl_logic;
        lsc_prog_incr_rti_c: in     vl_logic;
        lsc_prog_incr_enc_c: in     vl_logic;
        lsc_prog_incr_cmp_c: in     vl_logic;
        lsc_prog_incr_cne_c: in     vl_logic;
        lsc_vfy_incr_rti_c: in     vl_logic;
        lsc_prog_ctrl0_c: in     vl_logic;
        lsc_read_ctrl0_c: in     vl_logic;
        lsc_reset_crc_c : in     vl_logic;
        lsc_read_crc_c  : in     vl_logic;
        lsc_prog_sed_crc_c: in     vl_logic;
        lsc_read_sed_crc_c: in     vl_logic;
        lsc_prog_password_c: in     vl_logic;
        lsc_read_password_c: in     vl_logic;
        lsc_prog_cipher_key_c: in     vl_logic;
        lsc_read_cipher_key_c: in     vl_logic;
        lsc_prog_feature_c: in     vl_logic;
        lsc_read_feature_c: in     vl_logic;
        lsc_prog_feabits_c: in     vl_logic;
        lsc_read_feabits_c: in     vl_logic;
        lsc_prog_otps_c : in     vl_logic;
        lsc_read_otps_c : in     vl_logic;
        lsc_write_comp_dic_c: in     vl_logic;
        lsc_write_bus_addr_c: in     vl_logic;
        lsc_pcs_write_c : in     vl_logic;
        lsc_pcs_read_c  : in     vl_logic;
        lsc_ebr_write_c : in     vl_logic;
        lsc_ebr_read_c  : in     vl_logic;
        lsc_prog_incr_nv_c: in     vl_logic;
        lsc_read_incr_nv_c: in     vl_logic;
        lsc_init_addr_ufm_c: in     vl_logic;
        lsc_prog_tag_c  : in     vl_logic;
        lsc_erase_tag_c : in     vl_logic;
        lsc_read_tag_c  : in     vl_logic;
        lsc_chip_select_c: in     vl_logic;
        lsc_flow_through_c: in     vl_logic;
        lsc_jump_c      : in     vl_logic;
        nj_invalid_c    : in     vl_logic;
        sed_prog_incr_rti_cq: in     vl_logic;
        sed_prog_incr_cmp_cq: in     vl_logic;
        isc_nj_enabled  : in     vl_logic;
        isc_nj_disable_completing: in     vl_logic
    );
end njtag_logic;
