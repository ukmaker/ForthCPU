library verilog;
use verilog.vl_types.all;
entity sbnx4v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end sbnx4v1s;
