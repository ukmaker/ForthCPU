library verilog;
use verilog.vl_types.all;
entity CKHS_BUFX16 is
    port(
        z               : out    vl_logic;
        a               : in     vl_logic
    );
end CKHS_BUFX16;
