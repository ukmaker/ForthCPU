library verilog;
use verilog.vl_types.all;
entity dig_top is
    port(
        vssp            : in     vl_logic;
        vccp            : in     vl_logic;
        gpio_in         : in     vl_logic_vector(9 downto 0);
        gpio_out        : out    vl_logic_vector(9 downto 0);
        gpio_oeb        : out    vl_logic_vector(9 downto 0);
        gpio_pldn_en    : out    vl_logic_vector(9 downto 0);
        scl_in          : in     vl_logic;
        sda_in          : in     vl_logic;
        sda_out         : out    vl_logic;
        fsafeb          : in     vl_logic;
        wdat_in         : in     vl_logic;
        rdat_out        : out    vl_logic;
        rdat_oeb        : out    vl_logic;
        wrclk           : in     vl_logic;
        resetb_in_pin   : in     vl_logic;
        reset_in_b      : out    vl_logic;
        por_n           : in     vl_logic;
        por_off         : out    vl_logic;
        resetb_out_pin  : out    vl_logic;
        ascclk_oeb      : out    vl_logic;
        ascclk_out      : out    vl_logic;
        dtpo_en         : out    vl_logic;
        dtpi_en         : out    vl_logic;
        ana_rst_b       : out    vl_logic;
        rst_abg_b       : out    vl_logic;
        vmon_hc_en      : out    vl_logic_vector(1 downto 0);
        mfg_vmon_bypass : out    vl_logic;
        vmon_odd        : in     vl_logic;
        vmona           : in     vl_logic_vector(10 downto 1);
        vmonb           : in     vl_logic_vector(10 downto 1);
        vmon_cfg_drvmcbus: out    vl_logic;
        vmon_cfg_dataout: out    vl_logic_vector(7 downto 0);
        vmon_cfg_datain : in     vl_logic_vector(7 downto 0);
        vmon_ldsshdw    : out    vl_logic;
        vmon_ldshdwreg  : out    vl_logic;
        vmon_ldmshdw    : out    vl_logic;
        vmon_rdshdw     : out    vl_logic;
        mfg_vmon        : out    vl_logic;
        rst_clk_gen_b   : out    vl_logic;
        imon_hc_en      : out    vl_logic_vector(1 downto 0);
        imon_fcout      : in     vl_logic;
        imon_gf_a       : in     vl_logic;
        imon_gf_b       : in     vl_logic;
        imonhv_fcout    : in     vl_logic;
        imonhv_gf_a     : in     vl_logic;
        imonhv_gf_b     : in     vl_logic;
        cfg_imon        : out    vl_logic_vector(30 downto 0);
        mfg_imon        : out    vl_logic_vector(6 downto 0);
        hvout_data      : out    vl_logic_vector(4 downto 1);
        cfg_hvout       : out    vl_logic_vector(31 downto 0);
        safestate       : out    vl_logic;
        vdac_chan       : in     vl_logic_vector(2 downto 0);
        vdac_ready      : in     vl_logic;
        vdac_init       : in     vl_logic;
        vdacin          : out    vl_logic_vector(7 downto 0);
        vdac_resetb     : out    vl_logic;
        vdac_bpz        : out    vl_logic_vector(1 downto 0);
        vdac_trimoutenable: out    vl_logic_vector(3 downto 0);
        vdac_trim_dac   : out    vl_logic_vector(3 downto 0);
        mfg_vdac        : out    vl_logic_vector(4 downto 0);
        sync_sample     : in     vl_logic;
        tmon_betacomp   : in     vl_logic;
        tmon_modout     : in     vl_logic;
        tmon_demratio   : out    vl_logic_vector(15 downto 0);
        tmon_demout     : out    vl_logic;
        tmon_single_e   : out    vl_logic;
        tmon_chansel    : out    vl_logic_vector(2 downto 0);
        tmon_betabits   : out    vl_logic_vector(5 downto 0);
        tmon_beta_en    : out    vl_logic;
        tmon_beta_done  : out    vl_logic;
        tmon_adc_resetb : out    vl_logic;
        tmon_adc_clk    : out    vl_logic;
        tmon_porkchop   : out    vl_logic;
        mfg_tmon        : out    vl_logic_vector(7 downto 0);
        trim_tmon       : out    vl_logic;
        trim_se_deriv   : out    vl_logic;
        tmon_1a         : in     vl_logic;
        tmon_1b         : in     vl_logic;
        tmon_2a         : in     vl_logic;
        tmon_2b         : in     vl_logic;
        tmonint_1a      : in     vl_logic;
        tmonint_1b      : in     vl_logic;
        i2cdet_compout  : in     vl_logic;
        i2cdet_tapsel   : out    vl_logic_vector(2 downto 0);
        i2cdet_resetb   : out    vl_logic;
        i2cdet_clk      : out    vl_logic;
        mfg_i2cdet      : out    vl_logic;
        saradc_done     : in     vl_logic;
        mfg_sar_m_en    : out    vl_logic;
        mfg_sar_p_en    : out    vl_logic;
        saradc_atten    : out    vl_logic;
        saradc_socb     : out    vl_logic;
        saradc_data     : in     vl_logic_vector(9 downto 0);
        saradc_muxsel   : out    vl_logic_vector(3 downto 0);
        bg_caldone      : in     vl_logic;
        mfg_abg         : out    vl_logic_vector(12 downto 0);
        trim_bg_buff    : out    vl_logic_vector(27 downto 0);
        mfg_sp          : out    vl_logic_vector(3 downto 0);
        trim_sp_bg      : out    vl_logic_vector(4 downto 0);
        rst_osc_b       : out    vl_logic;
        rst_osc_tmr_b   : out    vl_logic;
        clk_loss_off    : out    vl_logic;
        wrclk_lost      : in     vl_logic;
        mclk            : out    vl_logic;
        mclkout         : in     vl_logic;
        trim_osc        : out    vl_logic_vector(3 downto 0);
        trim_osc_vref   : out    vl_logic_vector(2 downto 0);
        mfg_osc_vref    : out    vl_logic;
        mfg_en_dtpo     : out    vl_logic;
        mfg_en_dtpi     : out    vl_logic;
        mfg_en_atp1     : out    vl_logic;
        mfg_en_atp2     : out    vl_logic;
        mfg_en_matp1    : out    vl_logic;
        mfg_en_matp2    : out    vl_logic;
        mfg_vmon_enb    : out    vl_logic;
        mfg_dac_enb     : out    vl_logic;
        mfg_adc_enb     : out    vl_logic;
        mfg_abg_enb     : out    vl_logic;
        mfg_hvblk_dis   : out    vl_logic;
        dtpi            : in     vl_logic;
        cfgarray_dataout: out    vl_logic_vector(7 downto 0);
        volarray_dataout: out    vl_logic_vector(7 downto 0);
        mc_mcb_out      : out    vl_logic_vector(7 downto 0);
        i2c_dataout     : out    vl_logic_vector(7 downto 0);
        readid_out      : out    vl_logic_vector(7 downto 0);
        mfg_dataout     : out    vl_logic_vector(7 downto 0);
        cfgarray_datain : in     vl_logic_vector(7 downto 0);
        volarray_datain : in     vl_logic_vector(7 downto 0);
        mc_mcb_in       : in     vl_logic_vector(7 downto 0);
        i2c_datain      : in     vl_logic_vector(7 downto 0);
        mfg_datain      : in     vl_logic_vector(7 downto 0);
        cfgarray_dataout_oe: out    vl_logic;
        volarray_dataout_oe: out    vl_logic;
        mc_drvmcbus     : out    vl_logic;
        i2c_dataout_oe  : out    vl_logic;
        readid_drvmcbus : out    vl_logic;
        readmfg_drvmcbus: out    vl_logic;
        ee_flut_col_addr: out    vl_logic_vector(2 downto 0);
        ee_flut_row_addr: out    vl_logic_vector(3 downto 0);
        ee_twi_data     : out    vl_logic_vector(7 downto 0);
        ee_cfg_sel_array: out    vl_logic;
        ee_cfgtrim_drvmcbus: out    vl_logic;
        ee_cfgtrim_load_addrlat: out    vl_logic;
        ee_cfgtrim_load_datareg: out    vl_logic;
        ee_cfgtrim_sel_datareg: out    vl_logic;
        ee_data_enable  : out    vl_logic;
        ee_donebit_sel_array: out    vl_logic;
        ee_enable_erase : out    vl_logic;
        ee_enable_program: out    vl_logic;
        ee_faultlog_load_soft_datareg: out    vl_logic;
        ee_faultlog_sel_twi: out    vl_logic;
        ee_flut_drvmcbus: out    vl_logic;
        ee_flut_load_datareg: out    vl_logic;
        ee_flut_sel_array: out    vl_logic;
        ee_flut_sel_sdatareg: out    vl_logic;
        ee_i2cmsb_drvmcbus: out    vl_logic;
        ee_i2cmsb_load_datareg: out    vl_logic;
        ee_i2cmsb_sel_array: out    vl_logic;
        ee_mfg_cfgsel   : out    vl_logic;
        ee_mfg_dbg_iref : out    vl_logic;
        ee_mfg_dbg_vref : out    vl_logic;
        ee_mfg_donesel  : out    vl_logic;
        ee_mfg_faultsel : out    vl_logic;
        ee_mfg_i2csel   : out    vl_logic;
        ee_mfg_mcgforce : out    vl_logic;
        ee_mfg_mcgoe    : out    vl_logic;
        ee_mfg_progallrows: out    vl_logic;
        ee_mfg_progoddeve: out    vl_logic;
        ee_mfg_trimsel  : out    vl_logic;
        ee_mfg_vhien    : out    vl_logic;
        ee_mfg_vpp_pf   : out    vl_logic;
        ee_mfg_vppdiv   : out    vl_logic;
        ee_mfg_vppen    : out    vl_logic;
        ee_mfg_vppoe    : out    vl_logic;
        ee_vpptrim_erase: out    vl_logic_vector(4 downto 0);
        ee_vpptrim_program: out    vl_logic_vector(4 downto 0);
        ee_vbgtrim_reg  : out    vl_logic_vector(2 downto 0);
        ee_trim_sel_array: out    vl_logic;
        ee_slrtrim_reg  : out    vl_logic_vector(2 downto 0);
        ee_ibgtrim_reg  : out    vl_logic_vector(2 downto 0);
        ee_donebit      : in     vl_logic;
        ee_i2csa_done   : in     vl_logic;
        ee_i2csa        : in     vl_logic_vector(6 downto 3);
        ee_i2csa_lsb    : out    vl_logic_vector(2 downto 0)
    );
end dig_top;
