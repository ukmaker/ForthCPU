library verilog;
use verilog.vl_types.all;
entity asc_reno_mfg_array is
    generic(
        ASC_RENO        : integer := 1;
        ASC_VEGAS       : integer := 0;
        ASC_PROG_KEY_MSBYTE: integer := 229;
        ASC_PROG_KEY_LSBYTE: integer := 61;
        ASC_MFG_KEY_MSBYTE: integer := 156;
        ASC_MFG_KEY_LSBYTE: integer := 183;
        ASC_CFG_SIZE    : integer := 112;
        ASC_REG_WRALLRECFG_START: integer := 0;
        ASC_REG_CH1_PROFILE1_SETPOINT_LO: integer := 0;
        ASC_MSK_CH1_PROFILE1_SETPOINT_LO: integer := 255;
        ASC_REG_CH1_CH2_PROFILE1_SETPOINT_HI: integer := 1;
        ASC_MSK_CH1_CH2_PROFILE1_SETPOINT_HI: integer := 255;
        ASC_REG_CH2_PROFILE1_SETPOINT_LO: integer := 2;
        ASC_MSK_CH2_PROFILE1_SETPOINT_LO: integer := 255;
        ASC_REG_CH3_PROFILE1_SETPOINT_LO: integer := 3;
        ASC_MSK_CH3_PROFILE1_SETPOINT_LO: integer := 255;
        ASC_REG_CH3_CH4_PROFILE1_SETPOINT_HI: integer := 4;
        ASC_MSK_CH3_CH4_PROFILE1_SETPOINT_HI: integer := 255;
        ASC_REG_CH4_PROFILE1_SETPOINT_LO: integer := 5;
        ASC_MSK_CH4_PROFILE1_SETPOINT_LO: integer := 255;
        ASC_REG_CH1_PROFILE2_SETPOINT_LO: integer := 6;
        ASC_MSK_CH1_PROFILE2_SETPOINT_LO: integer := 255;
        ASC_REG_CH1_CH2_PROFILE2_SETPOINT_HI: integer := 7;
        ASC_MSK_CH1_CH2_PROFILE2_SETPOINT_HI: integer := 255;
        ASC_REG_CH2_PROFILE2_SETPOINT_LO: integer := 8;
        ASC_MSK_CH2_PROFILE2_SETPOINT_LO: integer := 255;
        ASC_REG_CH3_PROFILE2_SETPOINT_LO: integer := 9;
        ASC_MSK_CH3_PROFILE2_SETPOINT_LO: integer := 255;
        ASC_REG_CH3_CH4_PROFILE2_SETPOINT_HI: integer := 10;
        ASC_MSK_CH3_CH4_PROFILE2_SETPOINT_HI: integer := 255;
        ASC_REG_CH4_PROFILE2_SETPOINT_LO: integer := 11;
        ASC_MSK_CH4_PROFILE2_SETPOINT_LO: integer := 255;
        ASC_REG_CH1_PROFILE0_SETPOINT_LO: integer := 12;
        ASC_MSK_CH1_PROFILE0_SETPOINT_LO: integer := 255;
        ASC_REG_CH1_PROFILE0_SETPOINT_HI: integer := 13;
        ASC_MSK_CH1_PROFILE0_SETPOINT_HI: integer := 239;
        ASC_REG_CH2_PROFILE0_SETPOINT_LO: integer := 14;
        ASC_MSK_CH2_PROFILE0_SETPOINT_LO: integer := 255;
        ASC_REG_CH2_PROFILE0_SETPOINT_HI: integer := 15;
        ASC_MSK_CH2_PROFILE0_SETPOINT_HI: integer := 239;
        ASC_REG_CH3_PROFILE0_SETPOINT_LO: integer := 16;
        ASC_MSK_CH3_PROFILE0_SETPOINT_LO: integer := 255;
        ASC_REG_CH3_PROFILE0_SETPOINT_HI: integer := 17;
        ASC_MSK_CH3_PROFILE0_SETPOINT_HI: integer := 239;
        ASC_REG_CH4_PROFILE0_SETPOINT_LO: integer := 18;
        ASC_MSK_CH4_PROFILE0_SETPOINT_LO: integer := 255;
        ASC_REG_CH4_PROFILE0_SETPOINT_HI: integer := 19;
        ASC_MSK_CH4_PROFILE0_SETPOINT_HI: integer := 239;
        ASC_REG_CLT_CR  : integer := 20;
        ASC_MSK_CLT_CR  : integer := 3;
        ASC_REG_VDAC_CR0: integer := 21;
        ASC_MSK_VDAC_CR0: integer := 255;
        ASC_REG_VMON1_CR0: integer := 22;
        ASC_MSK_VMON1_CR0: integer := 255;
        ASC_REG_VMON1_CR1: integer := 23;
        ASC_MSK_VMON1_CR1: integer := 255;
        ASC_REG_VMON1_CR2: integer := 24;
        ASC_MSK_VMON1_CR2: integer := 255;
        ASC_REG_VMON2_CR0: integer := 25;
        ASC_MSK_VMON2_CR0: integer := 255;
        ASC_REG_VMON2_CR1: integer := 26;
        ASC_MSK_VMON2_CR1: integer := 255;
        ASC_REG_VMON2_CR2: integer := 27;
        ASC_MSK_VMON2_CR2: integer := 255;
        ASC_REG_VMON3_CR0: integer := 28;
        ASC_MSK_VMON3_CR0: integer := 255;
        ASC_REG_VMON3_CR1: integer := 29;
        ASC_MSK_VMON3_CR1: integer := 255;
        ASC_REG_VMON3_CR2: integer := 30;
        ASC_MSK_VMON3_CR2: integer := 255;
        ASC_REG_VMON4_CR0: integer := 31;
        ASC_MSK_VMON4_CR0: integer := 255;
        ASC_REG_VMON4_CR1: integer := 32;
        ASC_MSK_VMON4_CR1: integer := 255;
        ASC_REG_VMON4_CR2: integer := 33;
        ASC_MSK_VMON4_CR2: integer := 255;
        ASC_REG_VMON5_CR0: integer := 34;
        ASC_MSK_VMON5_CR0: integer := 255;
        ASC_REG_VMON5_CR1: integer := 35;
        ASC_MSK_VMON5_CR1: integer := 255;
        ASC_REG_VMON5_CR2: integer := 36;
        ASC_MSK_VMON5_CR2: integer := 255;
        ASC_REG_VMON6_CR0: integer := 37;
        ASC_MSK_VMON6_CR0: integer := 255;
        ASC_REG_VMON6_CR1: integer := 38;
        ASC_MSK_VMON6_CR1: integer := 255;
        ASC_REG_VMON6_CR2: integer := 39;
        ASC_MSK_VMON6_CR2: integer := 255;
        ASC_REG_VMON7_CR0: integer := 40;
        ASC_MSK_VMON7_CR0: integer := 255;
        ASC_REG_VMON7_CR1: integer := 41;
        ASC_MSK_VMON7_CR1: integer := 255;
        ASC_REG_VMON7_CR2: integer := 42;
        ASC_MSK_VMON7_CR2: integer := 255;
        ASC_REG_VMON8_CR0: integer := 43;
        ASC_MSK_VMON8_CR0: integer := 255;
        ASC_REG_VMON8_CR1: integer := 44;
        ASC_MSK_VMON8_CR1: integer := 255;
        ASC_REG_VMON8_CR2: integer := 45;
        ASC_MSK_VMON8_CR2: integer := 255;
        ASC_REG_VMON9_CR0: integer := 46;
        ASC_MSK_VMON9_CR0: integer := 255;
        ASC_REG_VMON9_CR1: integer := 47;
        ASC_MSK_VMON9_CR1: integer := 255;
        ASC_REG_VMON9_CR2: integer := 48;
        ASC_MSK_VMON9_CR2: integer := 255;
        ASC_REG_HVMON_CR0: integer := 49;
        ASC_MSK_HVMON_CR0: integer := 255;
        ASC_REG_HVMON_CR1: integer := 50;
        ASC_MSK_HVMON_CR1: integer := 255;
        ASC_REG_HVMON_CR2: integer := 51;
        ASC_MSK_HVMON_CR2: integer := 255;
        ASC_REG_IMON1_CR0: integer := 52;
        ASC_MSK_IMON1_CR0: integer := 255;
        ASC_REG_IMON1_CR1: integer := 53;
        ASC_MSK_IMON1_CR1: integer := 255;
        ASC_REG_HIMON1_CR0: integer := 54;
        ASC_MSK_HIMON1_CR0: integer := 251;
        ASC_REG_HIMON1_CR1: integer := 55;
        ASC_MSK_HIMON1_CR1: integer := 255;
        ASC_REG_TMON1_CR0: integer := 56;
        ASC_MSK_TMON1_CR0: integer := 255;
        ASC_REG_TMON1_CR1: integer := 57;
        ASC_MSK_TMON1_CR1: integer := 255;
        ASC_REG_TMON1_CR2: integer := 58;
        ASC_MSK_TMON1_CR2: integer := 255;
        ASC_REG_TMON1_CR3: integer := 59;
        ASC_MSK_TMON1_CR3: integer := 255;
        ASC_REG_TMON1_CR4: integer := 60;
        ASC_MSK_TMON1_CR4: integer := 255;
        ASC_REG_TMON1_CR5: integer := 61;
        ASC_MSK_TMON1_CR5: integer := 63;
        ASC_REG_TMON1_CR6: integer := 62;
        ASC_MSK_TMON1_CR6: integer := 255;
        ASC_REG_TMON1_CR7: integer := 63;
        ASC_MSK_TMON1_CR7: integer := 127;
        ASC_REG_TMON1_CR8: integer := 64;
        ASC_MSK_TMON1_CR8: integer := 127;
        ASC_REG_TMON2_CR0: integer := 65;
        ASC_MSK_TMON2_CR0: integer := 255;
        ASC_REG_TMON2_CR1: integer := 66;
        ASC_MSK_TMON2_CR1: integer := 255;
        ASC_REG_TMON2_CR2: integer := 67;
        ASC_MSK_TMON2_CR2: integer := 255;
        ASC_REG_TMON2_CR3: integer := 68;
        ASC_MSK_TMON2_CR3: integer := 255;
        ASC_REG_TMON2_CR4: integer := 69;
        ASC_MSK_TMON2_CR4: integer := 255;
        ASC_REG_TMON2_CR5: integer := 70;
        ASC_MSK_TMON2_CR5: integer := 63;
        ASC_REG_TMON2_CR6: integer := 71;
        ASC_MSK_TMON2_CR6: integer := 255;
        ASC_REG_TMON2_CR7: integer := 72;
        ASC_MSK_TMON2_CR7: integer := 127;
        ASC_REG_TMON2_CR8: integer := 73;
        ASC_MSK_TMON2_CR8: integer := 127;
        ASC_REG_TMONINT_CR0: integer := 74;
        ASC_MSK_TMONINT_CR0: integer := 255;
        ASC_REG_TMONINT_CR1: integer := 75;
        ASC_MSK_TMONINT_CR1: integer := 255;
        ASC_REG_TMONINT_CR2: integer := 76;
        ASC_MSK_TMONINT_CR2: integer := 255;
        ASC_REG_TMONINT_CR3: integer := 77;
        ASC_MSK_TMONINT_CR3: integer := 255;
        ASC_REG_TMONINT_CR4: integer := 78;
        ASC_MSK_TMONINT_CR4: integer := 255;
        ASC_REG_TMONINT_CR5: integer := 79;
        ASC_MSK_TMONINT_CR5: integer := 31;
        ASC_REG_TMONINT_CR6: integer := 80;
        ASC_MSK_TMONINT_CR6: integer := 255;
        ASC_REG_TMONINT_CR7: integer := 81;
        ASC_MSK_TMONINT_CR7: integer := 127;
        ASC_REG_TMONINT_CR8: integer := 82;
        ASC_MSK_TMONINT_CR8: integer := 127;
        ASC_REG_HVOUT1_CR0: integer := 83;
        ASC_MSK_HVOUT1_CR0: integer := 255;
        ASC_REG_HVOUT1_CR1: integer := 84;
        ASC_MSK_HVOUT1_CR1: integer := 239;
        ASC_REG_HVOUT2_CR0: integer := 85;
        ASC_MSK_HVOUT2_CR0: integer := 255;
        ASC_REG_HVOUT2_CR1: integer := 86;
        ASC_MSK_HVOUT2_CR1: integer := 239;
        ASC_REG_HVOUT3_CR0: integer := 87;
        ASC_MSK_HVOUT3_CR0: integer := 255;
        ASC_REG_HVOUT3_CR1: integer := 88;
        ASC_MSK_HVOUT3_CR1: integer := 239;
        ASC_REG_HVOUT4_CR0: integer := 89;
        ASC_MSK_HVOUT4_CR0: integer := 255;
        ASC_REG_HVOUT4_CR1: integer := 90;
        ASC_MSK_HVOUT4_CR1: integer := 239;
        ASC_REG_GCS_CR0 : integer := 91;
        ASC_MSK_GCS_CR0 : integer := 255;
        ASC_REG_GCS_CR1 : integer := 92;
        ASC_MSK_GCS_CR1 : integer := 255;
        ASC_REG_GCS_CR2 : integer := 93;
        ASC_MSK_GCS_CR2 : integer := 255;
        ASC_REG_GCS_CR3 : integer := 94;
        ASC_MSK_GCS_CR3 : integer := 63;
        ASC_REG_GCS_CR4 : integer := 95;
        ASC_MSK_GCS_CR4 : integer := 63;
        ASC_REG_GCS_CR5 : integer := 96;
        ASC_MSK_GCS_CR5 : integer := 127;
        ASC_REG_GPIO_SRC_SEL: integer := 97;
        ASC_MSK_GPIO_SRC_SEL: integer := 0;
        ASC_REG_GPIO_4_1_CR: integer := 98;
        ASC_MSK_GPIO_4_1_CR: integer := 85;
        ASC_REG_GPIO_8_5_CR: integer := 99;
        ASC_MSK_GPIO_8_5_CR: integer := 85;
        ASC_REG_GPIO_10_9_CR: integer := 100;
        ASC_MSK_GPIO_10_9_CR: integer := 5;
        ASC_REG_ASCCLK_DIS_CR: integer := 101;
        ASC_MSK_ASCCLK_DIS_CR: integer := 1;
        ASC_REG_WRITE_PROTECT_CR: integer := 102;
        ASC_MSK_WRITE_PROTECT_CR: integer := 3;
        ASC_REG_RSVD_CR0: integer := 103;
        ASC_MSK_RSVD_CR0: integer := 0;
        ASC_REG_RSVD_CR1: integer := 104;
        ASC_MSK_RSVD_CR1: integer := 0;
        ASC_REG_RSVD_CR2: integer := 105;
        ASC_MSK_RSVD_CR2: integer := 0;
        ASC_REG_RSVD_CR3: integer := 112;
        ASC_MSK_RSVD_CR3: integer := 0;
        ASC_REG_RSVD_CR4: integer := 107;
        ASC_MSK_RSVD_CR4: integer := 0;
        ASC_REG_RSVD_CR5: integer := 108;
        ASC_MSK_RSVD_CR5: integer := 0;
        ASC_REG_RSVD_CR6: integer := 109;
        ASC_MSK_RSVD_CR6: integer := 0;
        ASC_REG_RSVD_CR7: integer := 110;
        ASC_MSK_RSVD_CR7: integer := 0;
        ASC_REG_RSVD_CR8: integer := 111;
        ASC_MSK_RSVD_CR8: integer := 0;
        ASC_CSR_ADC_CONV_REQUEST: integer := 0;
        ASC_MSK_ADC_CONV_REQUEST: integer := 159;
        ASC_CSR_ADC_CONV_RESULT_LO: integer := 1;
        ASC_MSK_ADC_CONV_RESULT_LO: integer := 255;
        ASC_CSR_ADC_CONV_RESULT_HI: integer := 2;
        ASC_MSK_ADC_CONV_RESULT_HI: integer := 255;
        ASC_CSR_IMON_MAVG_CONTROL: integer := 3;
        ASC_MSK_IMON_MAVG_CONTROL: integer := 167;
        ASC_CSR_IMON_MAVG_SELECT: integer := 4;
        ASC_MSK_IMON_MAVG_SELECT: integer := 3;
        ASC_CSR_IMON_MAVG_RESULT_LO: integer := 5;
        ASC_MSK_IMON_MAVG_RESULT_LO: integer := 255;
        ASC_CSR_IMON_MAVG_RESULT_HI: integer := 6;
        ASC_MSK_IMON_MAVG_RESULT_HI: integer := 3;
        ASC_CSR_RDAT_MONITOR_CR: integer := 7;
        ASC_MSK_RDAT_MONITOR_CR: integer := 143;
        ASC_CSR_RDAT_MONITOR_DATA: integer := 8;
        ASC_MSK_RDAT_MONITOR_DATA: integer := 255;
        ASC_CSR_GCS_I2C_CTRL: integer := 112;
        ASC_MSK_GCS_I2C_CTRL: integer := 63;
        ASC_CSR_TMON_MEAS_CH0_HI_REG: integer := 128;
        ASC_MSK_TMON_MEAS_CH0_HI_REG: integer := 255;
        ASC_CSR_TMON_MEAS_CH0_LO_REG: integer := 129;
        ASC_MSK_TMON_MEAS_CH0_LO_REG: integer := 224;
        ASC_CSR_TMON_MEAS_CH1_HI_REG: integer := 130;
        ASC_MSK_TMON_MEAS_CH1_HI_REG: integer := 255;
        ASC_CSR_TMON_MEAS_CH1_LO_REG: integer := 131;
        ASC_MSK_TMON_MEAS_CH1_LO_REG: integer := 224;
        ASC_CSR_TMON_MEAS_CH2_HI_REG: integer := 132;
        ASC_MSK_TMON_MEAS_CH2_HI_REG: integer := 255;
        ASC_CSR_TMON_MEAS_CH2_LO_REG: integer := 133;
        ASC_MSK_TMON_MEAS_CH2_LO_REG: integer := 224;
        ASC_CSR_TMON_A_ALARM: integer := 134;
        ASC_MSK_TMON_A_ALARM: integer := 7;
        ASC_CSR_TMON_B_ALARM: integer := 135;
        ASC_MSK_TMON_B_ALARM: integer := 7;
        ASC_CSR_TMON_STATUS: integer := 136;
        ASC_MSK_TMON_STATUS: integer := 7;
        ASC_CSR_TMON_BETA_SAR: integer := 137;
        ASC_MSK_TMON_BETA_SAR: integer := 63;
        ASC_CSR_TMON_ANA_TEST: integer := 138;
        ASC_MSK_TMON_ANA_TEST: integer := 255;
        ASC_CSR_TMON_DIGFORANA_TEST: integer := 139;
        ASC_MSK_TMON_DIGFORANA_TEST: integer := 255;
        ASC_CSR_TMON_FILTER_DATA_LO: integer := 140;
        ASC_MSK_TMON_FILTER_DATA_LO: integer := 255;
        ASC_CSR_TMON_FILTER_DATA_HI: integer := 141;
        ASC_MSK_TMON_FILTER_DATA_HI: integer := 255;
        ASC_CSR_TMON_CTRL: integer := 142;
        ASC_MSK_TMON_CTRL: integer := 7;
        ASC_CSR_TMON_ALU_M_LO: integer := 143;
        ASC_MSK_TMON_ALU_M_LO: integer := 255;
        ASC_CSR_TMON_ALU_M_MLO: integer := 144;
        ASC_MSK_TMON_ALU_M_MLO: integer := 255;
        ASC_CSR_TMON_ALU_M_MHI: integer := 145;
        ASC_MSK_TMON_ALU_M_MHI: integer := 255;
        ASC_CSR_TMON_ALU_M_HI: integer := 146;
        ASC_MSK_TMON_ALU_M_HI: integer := 255;
        ASC_CSR_TMON_ALU_ACC_LO: integer := 147;
        ASC_MSK_TMON_ALU_ACC_LO: integer := 255;
        ASC_CSR_TMON_ALU_ACC_MLO: integer := 148;
        ASC_MSK_TMON_ALU_ACC_MLO: integer := 255;
        ASC_CSR_TMON_ALU_ACC_MHI: integer := 149;
        ASC_MSK_TMON_ALU_ACC_MHI: integer := 255;
        ASC_CSR_TMON_ALU_ACC_HI: integer := 150;
        ASC_MSK_TMON_ALU_ACC_HI: integer := 255;
        ASC_CSR_TMON_ALU_Q_LO: integer := 151;
        ASC_MSK_TMON_ALU_Q_LO: integer := 255;
        ASC_CSR_TMON_ALU_Q_MD: integer := 152;
        ASC_MSK_TMON_ALU_Q_MD: integer := 255;
        ASC_CSR_TMON_ALU_Q_HI: integer := 153;
        ASC_MSK_TMON_ALU_Q_HI: integer := 1;
        ASC_CSR_TMON_ALU_CMD: integer := 154;
        ASC_MSK_TMON_ALU_CMD: integer := 7;
        ASC_CSR_VALUE_VDAC1: integer := 160;
        ASC_MSK_VALUE_VDAC1: integer := 255;
        ASC_CSR_VALUE_VDAC2: integer := 161;
        ASC_MSK_VALUE_VDAC2: integer := 255;
        ASC_CSR_VALUE_VDAC3: integer := 162;
        ASC_MSK_VALUE_VDAC3: integer := 255;
        ASC_CSR_VALUE_VDAC4: integer := 163;
        ASC_MSK_VALUE_VDAC4: integer := 255;
        ASC_CSR_CLT_TST0: integer := 164;
        ASC_MSK_CLT_TST0: integer := 255;
        ASC_CSR_CLT_TST1: integer := 165;
        ASC_MSK_CLT_TST1: integer := 131;
        ASC_TRIM_BYTE_0 : integer := 0;
        ASC_TRIM_MSK_BYTE_0: integer := 255;
        ASC_TRIM_BYTE_1 : integer := 1;
        ASC_TRIM_MSK_BYTE_1: integer := 255;
        ASC_TRIM_BYTE_2 : integer := 2;
        ASC_TRIM_MSK_BYTE_2: integer := 255;
        ASC_TRIM_BYTE_3 : integer := 3;
        ASC_TRIM_MSK_BYTE_3: integer := 255;
        ASC_TRIM_BYTE_4 : integer := 4;
        ASC_TRIM_MSK_BYTE_4: integer := 255;
        ASC_TRIM_BYTE_5 : integer := 5;
        ASC_TRIM_MSK_BYTE_5: integer := 255;
        ASC_TRIM_BYTE_6 : integer := 6;
        ASC_TRIM_MSK_BYTE_6: integer := 1;
        ASC_TRIM_BYTE_7 : integer := 7;
        ASC_TRIM_MSK_BYTE_7: integer := 255;
        ASC_TRIM_BYTE_8 : integer := 8;
        ASC_TRIM_MSK_BYTE_8: integer := 239;
        ASC_TRIM_BYTE_9 : integer := 9;
        ASC_TRIM_MSK_BYTE_9: integer := 255;
        ASC_TRIM_BYTE_10: integer := 10;
        ASC_TRIM_MSK_BYTE_10: integer := 0;
        ASC_TRIM_BYTE_11: integer := 11;
        ASC_TRIM_MSK_BYTE_11: integer := 255;
        ASC_TRIM_BYTE_12: integer := 12;
        ASC_TRIM_MSK_BYTE_12: integer := 255;
        ASC_TRIM_BYTE_13: integer := 13;
        ASC_TRIM_MSK_BYTE_13: integer := 207;
        ASC_TRIM_BYTE_14: integer := 14;
        ASC_TRIM_MSK_BYTE_14: integer := 255;
        ASC_TRIM_BYTE_15: integer := 15;
        ASC_TRIM_MSK_BYTE_15: integer := 255;
        ASC_TRIM_BYTE_16: integer := 16;
        ASC_TRIM_MSK_BYTE_16: integer := 0;
        ASC_TRIM_BYTE_17: integer := 17;
        ASC_TRIM_MSK_BYTE_17: integer := 0;
        ASC_TRIM_BYTE_18: integer := 18;
        ASC_TRIM_MSK_BYTE_18: integer := 0;
        ASC_TRIM_BYTE_19: integer := 19;
        ASC_TRIM_MSK_BYTE_19: integer := 0;
        ASC_TRIM_BYTE_20: integer := 20;
        ASC_TRIM_MSK_BYTE_20: integer := 0;
        ASC_TRIM_BYTE_21: integer := 21;
        ASC_TRIM_MSK_BYTE_21: integer := 0;
        ASC_TRIM_BYTE_22: integer := 22;
        ASC_TRIM_MSK_BYTE_22: integer := 0;
        ASC_TRIM_BYTE_23: integer := 23;
        ASC_TRIM_MSK_BYTE_23: integer := 0;
        ASC_TRIM_BYTE_24: integer := 24;
        ASC_TRIM_MSK_BYTE_24: integer := 0;
        ASC_TRIM_BYTE_25: integer := 25;
        ASC_TRIM_MSK_BYTE_25: integer := 0;
        ASC_TRIM_BYTE_26: integer := 26;
        ASC_TRIM_MSK_BYTE_26: integer := 0;
        ASC_TRIM_BYTE_27: integer := 27;
        ASC_TRIM_MSK_BYTE_27: integer := 0;
        ASC_TRIM_BYTE_28: integer := 28;
        ASC_TRIM_MSK_BYTE_28: integer := 0;
        ASC_TRIM_BYTE_29: integer := 29;
        ASC_TRIM_MSK_BYTE_29: integer := 0;
        ASC_TRIM_BYTE_30: integer := 30;
        ASC_TRIM_MSK_BYTE_30: integer := 0;
        ASC_TRIM_BYTE_31: integer := 31;
        ASC_TRIM_MSK_BYTE_31: integer := 0;
        ASC_MFG_BYTE_0  : integer := 0;
        ASC_MFG_BYTE_1  : integer := 1;
        ASC_MFG_BYTE_2  : integer := 2;
        ASC_MFG_RST_BYTE_2: integer := 0;
        ASC_MFG_MSK_BYTE_2: integer := 255;
        ASC_MFG_BYTE_3  : integer := 3;
        ASC_MFG_RST_BYTE_3: integer := 0;
        ASC_MFG_MSK_BYTE_3: integer := 255;
        ASC_MFG_BYTE_4  : integer := 4;
        ASC_MFG_RST_BYTE_4: integer := 0;
        ASC_MFG_MSK_BYTE_4: integer := 255;
        ASC_MFG_BYTE_5  : integer := 5;
        ASC_MFG_RST_BYTE_5: integer := 0;
        ASC_MFG_MSK_BYTE_5: integer := 255;
        ASC_MFG_BYTE_6  : integer := 6;
        ASC_MFG_RST_BYTE_6: integer := 0;
        ASC_MFG_MSK_BYTE_6: integer := 255;
        ASC_MFG_BYTE_7  : integer := 7;
        ASC_MFG_RST_BYTE_7: integer := 0;
        ASC_MFG_MSK_BYTE_7: integer := 255;
        ASC_MFG_BYTE_8  : integer := 8;
        ASC_MFG_RST_BYTE_8: integer := 0;
        ASC_MFG_MSK_BYTE_8: integer := 255;
        ASC_MFG_BYTE_9  : integer := 9;
        ASC_MFG_RST_BYTE_9: integer := 0;
        ASC_MFG_MSK_BYTE_9: integer := 255;
        ASC_MFG_BYTE_10 : integer := 10;
        ASC_MFG_RST_BYTE_10: integer := 0;
        ASC_MFG_MSK_BYTE_10: integer := 255;
        ASC_MFG_BYTE_11 : integer := 11;
        ASC_MFG_RST_BYTE_11: integer := 0;
        ASC_MFG_MSK_BYTE_11: integer := 255;
        ASC_MFG_BYTE_12 : integer := 12;
        ASC_MFG_RST_BYTE_12: integer := 0;
        ASC_MFG_MSK_BYTE_12: integer := 247;
        ASC_MFG_BYTE_13 : integer := 13;
        ASC_MFG_RST_BYTE_13: integer := 0;
        ASC_MFG_MSK_BYTE_13: integer := 255
    );
    port(
        mfgbus_ld_addr_latch: in     vl_logic;
        mfgbus_ld_master_data_latch: in     vl_logic;
        mfgbus_datain   : in     vl_logic_vector(7 downto 0);
        mfgbus_dataout  : out    vl_logic_vector(7 downto 0);
        mfgbus_resetn   : in     vl_logic;
        mfgbus_clock    : in     vl_logic;
        mfg_array_mfg_mode: out    vl_logic;
        mfg_array_mcgoe : out    vl_logic;
        mfg_array_mcgforce: out    vl_logic;
        mfg_array_cfgsel: out    vl_logic;
        mfg_array_trimsel: out    vl_logic;
        mfg_array_i2csel: out    vl_logic;
        mfg_array_faultsel: out    vl_logic;
        mfg_array_donesel: out    vl_logic;
        mfg_array_vppoe : out    vl_logic;
        mfg_array_vppen : out    vl_logic;
        mfg_array_vppdiv: out    vl_logic;
        mfg_array_poroff: out    vl_logic;
        mfg_array_vhien : out    vl_logic;
        mfg_array_clttst_en: out    vl_logic;
        mfg_array_int2  : out    vl_logic;
        mfg_array_int1  : out    vl_logic;
        mfg_array_int0  : out    vl_logic;
        mfg_array_hvblank_dis: out    vl_logic;
        mfg_array_vpp_pf: out    vl_logic;
        mfg_array_vdac_en: out    vl_logic;
        mfg_array_vdac4 : out    vl_logic;
        mfg_array_vdac3 : out    vl_logic;
        mfg_array_vdac2 : out    vl_logic;
        mfg_array_vdac1 : out    vl_logic;
        mfg_array_i2caddr_en: out    vl_logic;
        mfg_array_dbg_vref: out    vl_logic;
        mfg_array_dbg_iref: out    vl_logic;
        mfg_array_tmonclk_dis: out    vl_logic;
        mfg_array_vmon_enb: out    vl_logic;
        mfg_array_adc_enb: out    vl_logic;
        mfg_array_dac_enb: out    vl_logic;
        mfg_array_abg_enb: out    vl_logic;
        mfg_array_test_clk_en: out    vl_logic;
        mfg_array_osc_vref: out    vl_logic;
        mfg_array_tmon_tst_en: out    vl_logic;
        mfg_array_sp_mfg_3: out    vl_logic;
        mfg_array_sp_mfg_2: out    vl_logic;
        mfg_array_sp_mfg_1: out    vl_logic;
        mfg_array_sp_mfg_0: out    vl_logic;
        mfg_array_vmon_test: out    vl_logic;
        mfg_array_vmon_bypass: out    vl_logic;
        mfg_array_fc_enb: out    vl_logic;
        mfg_array_sc_enb: out    vl_logic;
        mfg_array_imhv_atp_en: out    vl_logic;
        mfg_array_imon_atp_en: out    vl_logic;
        mfg_array_mfgvcm_drop: out    vl_logic;
        mfg_array_pga_enb: out    vl_logic;
        mfg_array_mfg_pga_chk: out    vl_logic;
        mfg_xorbus_rdat_enable: out    vl_logic;
        mfg_array_vtc_4 : out    vl_logic;
        mfg_array_vtc_3 : out    vl_logic;
        mfg_array_vtc_2 : out    vl_logic;
        mfg_array_vtc_1 : out    vl_logic;
        mfg_array_vtc_0 : out    vl_logic;
        mfg_array_timer_tst_en: out    vl_logic;
        mfg_array_buf_cref_tst: out    vl_logic;
        mfg_array_buf_vdac_tst: out    vl_logic;
        mfg_array_buf_tmon_tst: out    vl_logic;
        mfg_array_a2d_test_vip_en: out    vl_logic;
        mfg_array_a2d_test_vim_en: out    vl_logic;
        mfg_array_abias_test_en: out    vl_logic;
        mfg_array_abgtreg_2: out    vl_logic;
        mfg_array_abgtreg_1: out    vl_logic;
        mfg_array_abgtreg_0: out    vl_logic;
        mfg_array_clklossdetect_dis: out    vl_logic;
        mfg_array_atp1_en: out    vl_logic;
        mfg_array_atp2_en: out    vl_logic;
        mfg_array_matp1_en: out    vl_logic;
        mfg_array_matp2_en: out    vl_logic;
        mfg_array_dtpi_en: out    vl_logic;
        mfg_array_dtpo_en: out    vl_logic;
        mfg_array_twi_crcpad_dis: out    vl_logic;
        mfg_array_twi_loopback_en: out    vl_logic;
        mfg_array_anarst_dis: out    vl_logic;
        mfg_array_abgrst_dis: out    vl_logic;
        mfg_array_i2caddr_vdac_rst_dis: out    vl_logic;
        mfg_array_oscresetb_en: out    vl_logic;
        mfg_array_abgcu_tst_en: out    vl_logic;
        mfg_array_clk_sync_en: out    vl_logic;
        mfg_array_progallrows: out    vl_logic;
        mfg_array_progoddeve: out    vl_logic;
        mfg_array_vdac_reset: out    vl_logic;
        mfg_array_mfg_en_dtpi: out    vl_logic;
        mfg_array_mfg_en_dtpo: out    vl_logic;
        mfg_array_abg_reset: out    vl_logic;
        mfg_vdac_input_en: out    vl_logic;
        mfg_vdac_mfg_bpz: out    vl_logic_vector(1 downto 0);
        mfg_vdac_mfg_data: out    vl_logic_vector(7 downto 0)
    );
end asc_reno_mfg_array;
