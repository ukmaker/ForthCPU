library verilog;
use verilog.vl_types.all;
entity cfg_qual is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 1
    );
    port(
        jump_exec       : out    vl_logic;
        chip_select_exec: out    vl_logic;
        flow_through_exec: out    vl_logic;
        bypass_exec     : out    vl_logic;
        isc_data_shift_iqual: out    vl_logic;
        lsc_prog_incr_rti_iqual: out    vl_logic;
        lsc_prog_incr_enc_iqual: out    vl_logic;
        lsc_prog_incr_cmp_iqual: out    vl_logic;
        lsc_prog_incr_cne_iqual: out    vl_logic;
        isc_data_shift_cqual: out    vl_logic;
        lsc_prog_incr_rti_cqual: out    vl_logic;
        lsc_prog_incr_enc_cqual: out    vl_logic;
        lsc_prog_incr_cmp_cqual: out    vl_logic;
        lsc_prog_incr_cne_cqual: out    vl_logic;
        verify_id_qual  : out    vl_logic;
        read_temp_qual  : out    vl_logic;
        lsc_device_ctrl_qual: out    vl_logic;
        lsc_shift_password_qual: out    vl_logic;
        lsc_bitstream_burst_qual: out    vl_logic;
        lsc_read_pes_qual: out    vl_logic;
        sf_address_shift_qual: out    vl_logic;
        lsc_prog_ctrl0_qual: out    vl_logic;
        lsc_read_ctrl0_qual: out    vl_logic;
        lsc_reset_crc_qual: out    vl_logic;
        lsc_read_crc_qual: out    vl_logic;
        lsc_write_comp_dic_qual: out    vl_logic;
        lsc_read_comp_dic_qual: out    vl_logic;
        sed_init_addr_qual: out    vl_logic;
        sed_write_addr_qual: out    vl_logic;
        sed_read_incr_qual: out    vl_logic;
        sed_prog_sed_crc_qual: out    vl_logic;
        sed_prog_ctrl0_qual: out    vl_logic;
        sed_write_comp_dic_qual: out    vl_logic;
        sf_prog_ucode_qual: out    vl_logic;
        sf_program_qual : out    vl_logic;
        sf_read_qual    : out    vl_logic;
        sf_erase_qual   : out    vl_logic;
        sf_prog_done_qual: out    vl_logic;
        sf_erase_done_qual: out    vl_logic;
        sf_prog_sec_qual: out    vl_logic;
        sf_init_addr_qual: out    vl_logic;
        sf_write_addr_qual: out    vl_logic;
        sf_prog_incr_rti_qual: out    vl_logic;
        sf_prog_incr_enc_qual: out    vl_logic;
        sf_prog_incr_cmp_qual: out    vl_logic;
        sf_prog_incr_cne_qual: out    vl_logic;
        sf_vfy_incr_rti_qual: out    vl_logic;
        sf_prog_sed_crc_qual: out    vl_logic;
        sf_read_sed_crc_qual: out    vl_logic;
        sf_write_bus_addr_qual: out    vl_logic;
        sf_pcs_write_qual: out    vl_logic;
        sf_pcs_read_qual: out    vl_logic;
        sf_ebr_write_qual: out    vl_logic;
        sf_ebr_read_qual: out    vl_logic;
        sf_prog_std_all : out    vl_logic;
        sf_prog_enc_all : out    vl_logic;
        fl_prog_ucode_qual: out    vl_logic;
        fl_erase_qual   : out    vl_logic;
        fl_prog_done_qual: out    vl_logic;
        fl_prog_sec_qual: out    vl_logic;
        fl_prog_secplus_qual: out    vl_logic;
        fl_init_addr_qual: out    vl_logic;
        fl_write_addr_qual: out    vl_logic;
        fl_prog_incr_nv_qual: out    vl_logic;
        fl_read_incr_nv_qual: out    vl_logic;
        fl_prog_password_qual: out    vl_logic;
        fl_prog_cipher_key_qual: out    vl_logic;
        fl_prog_feature_qual: out    vl_logic;
        fl_prog_feabits_qual: out    vl_logic;
        fl_prog_otps_qual: out    vl_logic;
        fl_init_addr_ufm_qual: out    vl_logic;
        fl_prog_tag_qual: out    vl_logic;
        fl_erase_tag_qual: out    vl_logic;
        fl_read_tag_qual: out    vl_logic;
        fl_prog_pes_qual: out    vl_logic;
        fl_prog_mes_qual: out    vl_logic;
        fl_prog_hes_qual: out    vl_logic;
        fl_prog_trim_qual: out    vl_logic;
        fl_read_hes_qual: out    vl_logic;
        fl_mtest_qual   : out    vl_logic;
        ef_init_addr_qual: out    vl_logic;
        ef_write_addr_qual: out    vl_logic;
        ef_prog_password_qual: out    vl_logic;
        ef_prog_cipher_key_qual: out    vl_logic;
        ef_prog_feature_qual: out    vl_logic;
        ef_prog_feabits_qual: out    vl_logic;
        ef_prog_otps_qual: out    vl_logic;
        ef_prog_pes_qual: out    vl_logic;
        ef_prog_mes_qual: out    vl_logic;
        ef_prog_hes_qual: out    vl_logic;
        ef_prog_trim_qual: out    vl_logic;
        ef_read_hes_qual: out    vl_logic;
        ef_mtest_qual   : out    vl_logic;
        isc_prog_done_qual: out    vl_logic;
        isc_prog_sec_qual: out    vl_logic;
        isc_prog_secplus_qual: out    vl_logic;
        lsc_prog_password_qual: out    vl_logic;
        lsc_prog_cipher_key_qual: out    vl_logic;
        lsc_prog_feature_qual: out    vl_logic;
        lsc_prog_feabits_qual: out    vl_logic;
        lsc_prog_otps_qual: out    vl_logic;
        lsc_prog_trim_qual: out    vl_logic;
        lsc_prog_pes_qual: out    vl_logic;
        lsc_prog_mes_qual: out    vl_logic;
        lsc_read_password_qual: out    vl_logic;
        lsc_read_cipher_key_qual: out    vl_logic;
        lsc_read_feature_qual: out    vl_logic;
        lsc_read_feabits_qual: out    vl_logic;
        lsc_read_otps_qual: out    vl_logic;
        lsc_read_trim_qual: out    vl_logic;
        lsc_read_mes_qual: out    vl_logic;
        mfg_mdata_qual  : out    vl_logic;
        mfg_mtrim_qual  : out    vl_logic;
        cmd_read_exec_buf: out    vl_logic;
        cmd_read_cfg_reg: out    vl_logic;
        cmd_prog_cfg_reg: out    vl_logic;
        bse_prog_incr_cqual: out    vl_logic;
        lsc_i2ci_crbr_wt_qual: out    vl_logic;
        lsc_i2ci_txdr_wt_qual: out    vl_logic;
        lsc_i2ci_rxdr_rd_qual: out    vl_logic;
        lsc_i2ci_sr_rd_qual: out    vl_logic;
        lsc_read_i2c_qual: out    vl_logic;
        pwd_mismatch_all: in     vl_logic;
        sd_key_lock     : in     vl_logic;
        sd_dec_only     : in     vl_logic;
        read_sram_dis   : in     vl_logic;
        write_sram_dis  : in     vl_logic;
        erase_sram_dis  : in     vl_logic;
        read_flfea_dis  : in     vl_logic;
        write_flfea_dis : in     vl_logic;
        erase_flfea_dis : in     vl_logic;
        read_otps_dis   : in     vl_logic;
        write_otps_dis  : in     vl_logic;
        read_flcfg_dis  : in     vl_logic;
        write_flcfg_dis : in     vl_logic;
        erase_flcfg_dis : in     vl_logic;
        read_flufm_dis  : in     vl_logic;
        write_flufm_dis : in     vl_logic;
        erase_flufm_dis : in     vl_logic;
        read_efuse_dis  : in     vl_logic;
        write_efuse_dis : in     vl_logic;
        njbse_rxdec     : in     vl_logic;
        p_mspi_all      : in     vl_logic;
        isc_exec_d      : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        mfg_margin_en   : in     vl_logic;
        cfg_sed_en      : in     vl_logic;
        dev_sdm_inp     : in     vl_logic;
        fl_row_sec      : in     vl_logic_vector(1 downto 0);
        isc_data_shift_iq: in     vl_logic;
        isc_addr_shift_iq: in     vl_logic;
        verify_id_iq    : in     vl_logic;
        read_temp_iq    : in     vl_logic;
        lsc_device_ctrl_iq: in     vl_logic;
        lsc_shift_password_iq: in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic;
        lsc_i2ci_crbr_wt_iq: in     vl_logic;
        lsc_i2ci_txdr_wt_iq: in     vl_logic;
        lsc_i2ci_rxdr_rd_iq: in     vl_logic;
        lsc_i2ci_sr_rd_iq: in     vl_logic;
        lsc_read_pes_mq : in     vl_logic;
        lsc_prog_ctrl0_iq: in     vl_logic;
        lsc_read_ctrl0_iq: in     vl_logic;
        lsc_reset_crc_iq: in     vl_logic;
        lsc_read_crc_iq : in     vl_logic;
        lsc_write_comp_dic_iq: in     vl_logic;
        lsc_read_comp_dic_mq: in     vl_logic;
        sf_prog_ucode_iq: in     vl_logic;
        sf_program_iq   : in     vl_logic;
        sf_read_iq      : in     vl_logic;
        sf_erase_iq     : in     vl_logic;
        sf_prog_done_iq : in     vl_logic;
        sf_erase_done_iq: in     vl_logic;
        sf_prog_sec_iq  : in     vl_logic;
        sf_init_addr_iq : in     vl_logic;
        sf_write_addr_iq: in     vl_logic;
        sf_prog_incr_rti_iq: in     vl_logic;
        sf_prog_incr_enc_iq: in     vl_logic;
        sf_prog_incr_cmp_iq: in     vl_logic;
        sf_prog_incr_cne_iq: in     vl_logic;
        sf_vfy_incr_rti_iq: in     vl_logic;
        sf_prog_sed_crc_iq: in     vl_logic;
        sf_read_sed_crc_iq: in     vl_logic;
        sf_write_bus_addr_iq: in     vl_logic;
        sf_pcs_write_iq : in     vl_logic;
        sf_pcs_read_iq  : in     vl_logic;
        sf_ebr_write_iq : in     vl_logic;
        sf_ebr_read_iq  : in     vl_logic;
        fl_prog_ucode_iq: in     vl_logic;
        fl_erase_iq     : in     vl_logic;
        fl_prog_done_iq : in     vl_logic;
        fl_prog_sec_iq  : in     vl_logic;
        fl_prog_secplus_iq: in     vl_logic;
        fl_init_addr_iq : in     vl_logic;
        fl_write_addr_iq: in     vl_logic;
        fl_prog_incr_nv_iq: in     vl_logic;
        fl_read_incr_nv_iq: in     vl_logic;
        fl_prog_password_iq: in     vl_logic;
        fl_read_password_iq: in     vl_logic;
        fl_prog_cipher_key_iq: in     vl_logic;
        fl_read_cipher_key_iq: in     vl_logic;
        fl_prog_feature_iq: in     vl_logic;
        fl_read_feature_iq: in     vl_logic;
        fl_prog_feabits_iq: in     vl_logic;
        fl_read_feabits_iq: in     vl_logic;
        fl_prog_otps_iq : in     vl_logic;
        fl_read_otps_iq : in     vl_logic;
        fl_init_addr_ufm_iq: in     vl_logic;
        fl_prog_tag_iq  : in     vl_logic;
        fl_erase_tag_iq : in     vl_logic;
        fl_read_tag_iq  : in     vl_logic;
        fl_prog_pes_mq  : in     vl_logic;
        fl_prog_trim_mq : in     vl_logic;
        fl_prog_mes_mq  : in     vl_logic;
        fl_prog_hes_mq  : in     vl_logic;
        fl_read_trim_mq : in     vl_logic;
        fl_read_mes_mq  : in     vl_logic;
        fl_read_hes_mq  : in     vl_logic;
        ef_init_addr_iq : in     vl_logic;
        ef_write_addr_iq: in     vl_logic;
        ef_prog_password_iq: in     vl_logic;
        ef_read_password_iq: in     vl_logic;
        ef_prog_cipher_key_iq: in     vl_logic;
        ef_read_cipher_key_iq: in     vl_logic;
        ef_prog_feature_iq: in     vl_logic;
        ef_read_feature_iq: in     vl_logic;
        ef_prog_feabits_iq: in     vl_logic;
        ef_read_feabits_iq: in     vl_logic;
        ef_prog_otps_iq : in     vl_logic;
        ef_read_otps_iq : in     vl_logic;
        ef_prog_pes_mq  : in     vl_logic;
        ef_prog_trim_mq : in     vl_logic;
        ef_prog_mes_mq  : in     vl_logic;
        ef_prog_hes_mq  : in     vl_logic;
        ef_read_trim_mq : in     vl_logic;
        ef_read_mes_mq  : in     vl_logic;
        ef_read_hes_mq  : in     vl_logic;
        mfg_mtest_mq    : in     vl_logic;
        mfg_mtrim_mq    : in     vl_logic;
        mfg_mdata_mq    : in     vl_logic;
        isc_data_shift_cq: in     vl_logic;
        isc_addr_shift_cq: in     vl_logic;
        verify_id_cq    : in     vl_logic;
        read_temp_cq    : in     vl_logic;
        lsc_device_ctrl_cq: in     vl_logic;
        lsc_shift_password_cq: in     vl_logic;
        lsc_bitstream_burst_cq: in     vl_logic;
        lsc_read_pes_cq : in     vl_logic;
        lsc_prog_ctrl0_cq: in     vl_logic;
        lsc_read_ctrl0_cq: in     vl_logic;
        lsc_reset_crc_cq: in     vl_logic;
        lsc_read_crc_cq : in     vl_logic;
        lsc_write_comp_dic_cq: in     vl_logic;
        sf_prog_ucode_cq: in     vl_logic;
        sf_program_cq   : in     vl_logic;
        sf_read_cq      : in     vl_logic;
        sf_erase_cq     : in     vl_logic;
        sf_prog_done_cq : in     vl_logic;
        sf_erase_done_cq: in     vl_logic;
        sf_prog_sec_cq  : in     vl_logic;
        sf_init_addr_cq : in     vl_logic;
        sf_write_addr_cq: in     vl_logic;
        sf_prog_incr_rti_cq: in     vl_logic;
        sf_prog_incr_enc_cq: in     vl_logic;
        sf_prog_incr_cmp_cq: in     vl_logic;
        sf_prog_incr_cne_cq: in     vl_logic;
        sf_vfy_incr_rti_cq: in     vl_logic;
        sf_prog_sed_crc_cq: in     vl_logic;
        sf_read_sed_crc_cq: in     vl_logic;
        sf_write_bus_addr_cq: in     vl_logic;
        sf_pcs_write_cq : in     vl_logic;
        sf_pcs_read_cq  : in     vl_logic;
        sf_ebr_write_cq : in     vl_logic;
        sf_ebr_read_cq  : in     vl_logic;
        fl_prog_ucode_cq: in     vl_logic;
        fl_erase_cq     : in     vl_logic;
        fl_prog_done_cq : in     vl_logic;
        fl_prog_sec_cq  : in     vl_logic;
        fl_prog_secplus_cq: in     vl_logic;
        fl_init_addr_cq : in     vl_logic;
        fl_write_addr_cq: in     vl_logic;
        fl_prog_incr_nv_cq: in     vl_logic;
        fl_read_incr_nv_cq: in     vl_logic;
        fl_prog_password_cq: in     vl_logic;
        fl_read_password_cq: in     vl_logic;
        fl_prog_cipher_key_cq: in     vl_logic;
        fl_read_cipher_key_cq: in     vl_logic;
        fl_prog_feature_cq: in     vl_logic;
        fl_read_feature_cq: in     vl_logic;
        fl_prog_feabits_cq: in     vl_logic;
        fl_read_feabits_cq: in     vl_logic;
        fl_prog_otps_cq : in     vl_logic;
        fl_read_otps_cq : in     vl_logic;
        fl_init_addr_ufm_cq: in     vl_logic;
        fl_prog_tag_cq  : in     vl_logic;
        fl_erase_tag_cq : in     vl_logic;
        fl_read_tag_cq  : in     vl_logic;
        ef_init_addr_cq : in     vl_logic;
        ef_write_addr_cq: in     vl_logic;
        ef_prog_password_cq: in     vl_logic;
        ef_read_password_cq: in     vl_logic;
        ef_prog_cipher_key_cq: in     vl_logic;
        ef_read_cipher_key_cq: in     vl_logic;
        ef_prog_feature_cq: in     vl_logic;
        ef_read_feature_cq: in     vl_logic;
        ef_prog_feabits_cq: in     vl_logic;
        ef_read_feabits_cq: in     vl_logic;
        ef_prog_otps_cq : in     vl_logic;
        ef_read_otps_cq : in     vl_logic;
        lsc_jump_cq     : in     vl_logic;
        lsc_chip_select_cq: in     vl_logic;
        lsc_flow_through_cq: in     vl_logic;
        bypass_cq       : in     vl_logic;
        sed_init_addr_cq: in     vl_logic;
        sed_write_addr_cq: in     vl_logic;
        sed_prog_incr_rti_cq: in     vl_logic;
        sed_prog_incr_cmp_cq: in     vl_logic;
        sed_prog_sed_crc_cq: in     vl_logic;
        sed_prog_ctrl0_cq: in     vl_logic;
        sed_write_comp_dic_cq: in     vl_logic;
        lsc_i2ci_crbr_wt_cq: in     vl_logic;
        lsc_i2ci_txdr_wt_cq: in     vl_logic;
        lsc_i2ci_rxdr_rd_cq: in     vl_logic;
        lsc_i2ci_sr_rd_cq: in     vl_logic
    );
end cfg_qual;
