library verilog;
use verilog.vl_types.all;
entity instruction is
    generic(
        ASC_I2C_INSTR_TRISTPAD: integer := 131;
        ASC_I2C_INSTR_LDRECFG: integer := 53;
        ASC_I2C_INSTR_SAFESTATE: integer := 130;
        ASC_I2C_INSTR_USERLOGICRST: integer := 129;
        ASC_I2C_INSTR_USERMODE: integer := 5;
        ASC_I2C_INSTR_LDSHDW: integer := 40;
        ASC_I2C_INSTR_BEUSER: integer := 6;
        ASC_I2C_INSTR_ERASEDONE: integer := 38;
        ASC_I2C_INSTR_PROGDONE: integer := 39;
        ASC_I2C_INSTR_ERASEI2CSA: integer := 17;
        ASC_I2C_INSTR_PROGI2CSA: integer := 20;
        ASC_I2C_INSTR_BECFG: integer := 33;
        ASC_I2C_INSTR_PROGCFG: integer := 36;
        ASC_I2C_INSTR_LDTRIMSHDW: integer := 149;
        ASC_I2C_INSTR_ERASEFAULT: integer := 113;
        ASC_I2C_INSTR_ERASEUSERTAG: integer := 97;
        ASC_I2C_INSTR_PROGUSERTAG: integer := 100;
        ASC_I2C_INSTR_BEALL: integer := 134;
        ASC_I2C_INSTR_PROGTRIM: integer := 147;
        ASC_I2C_INSTR_RDSHDW: integer := 51;
        ASC_I2C_INSTR_RDALLSHDW: integer := 52;
        ASC_I2C_INSTR_VERCFG: integer := 37;
        ASC_I2C_INSTR_VERUSERTAG: integer := 101;
        ASC_I2C_INSTR_RDSTATUS: integer := 3;
        ASC_I2C_INSTR_READI2CSA: integer := 19;
        ASC_I2C_INSTR_VERI2CSA: integer := 21;
        ASC_I2C_INSTR_RDTRIMSHDW: integer := 151;
        ASC_I2C_INSTR_RDFAULTEN: integer := 116;
        ASC_I2C_INSTR_RDID: integer := 2;
        ASC_I2C_INSTR_READCFG: integer := 35;
        ASC_I2C_INSTR_RDCFGCRC: integer := 55;
        ASC_I2C_INSTR_RDSOFTFAULT: integer := 115;
        ASC_I2C_INSTR_VERFAULT: integer := 117;
        ASC_I2C_INSTR_RDALLFAULT: integer := 118;
        ASC_I2C_INSTR_READUSERTAG: integer := 99;
        ASC_I2C_INSTR_READMFG: integer := 133;
        ASC_I2C_INSTR_READTRIM: integer := 146;
        ASC_I2C_INSTR_VERTRIM: integer := 148;
        ASC_I2C_INSTR_WRITECFG: integer := 34;
        ASC_I2C_INSTR_WRRECFG: integer := 49;
        ASC_I2C_INSTR_WRRECFGMASK: integer := 50;
        ASC_I2C_INSTR_WRALLRECFG: integer := 54;
        ASC_I2C_INSTR_WRRDVID1: integer := 65;
        ASC_I2C_INSTR_WRRDVID2: integer := 66;
        ASC_I2C_INSTR_WRRDVID3: integer := 67;
        ASC_I2C_INSTR_WRRDVID4: integer := 68;
        ASC_I2C_INSTR_WRRDVID5: integer := 69;
        ASC_I2C_INSTR_WRRDVID6: integer := 70;
        ASC_I2C_INSTR_WRRDVID7: integer := 71;
        ASC_I2C_INSTR_WRRDVID8: integer := 72;
        ASC_I2C_INSTR_WRITEUSERTAG: integer := 98;
        ASC_I2C_INSTR_WRITEMFG: integer := 132;
        ASC_I2C_INSTR_WRITETRIM: integer := 145;
        ASC_I2C_INSTR_ENPROG: integer := 4;
        ASC_I2C_INSTR_WRITEI2CSA: integer := 18;
        ASC_I2C_INSTR_WRTRIMSHDW: integer := 150;
        ASC_I2C_INSTR_TSTNRTHKEEPR: integer := 135;
        ASC_I2C_INSTR_WRMEASCTRL: integer := 81;
        ASC_I2C_INSTR_RDMEASRESULT: integer := 82;
        ASC_I2C_INSTR_NOOP: integer := 1
    );
    port(
        tristpad_iflg   : out    vl_logic;
        usermode_iflg   : out    vl_logic;
        ldshdw_iflg     : out    vl_logic;
        beuser_iflg     : out    vl_logic;
        erasedone_iflg  : out    vl_logic;
        progdone_iflg   : out    vl_logic;
        bei2csa_iflg    : out    vl_logic;
        progi2csa_iflg  : out    vl_logic;
        becfg_iflg      : out    vl_logic;
        progcfg_iflg    : out    vl_logic;
        eraseflut_iflg  : out    vl_logic;
        progusertag_iflg: out    vl_logic;
        eraseall_iflg   : out    vl_logic;
        progtrim_iflg   : out    vl_logic;
        rdshdw_iflg     : out    vl_logic;
        rdallshdw_iflg  : out    vl_logic;
        vercfg_iflg     : out    vl_logic;
        readstat_iflg   : out    vl_logic;
        rdi2csa_iflg    : out    vl_logic;
        veri2csa_iflg   : out    vl_logic;
        readid_iflg     : out    vl_logic;
        readcfg_iflg    : out    vl_logic;
        rdcfgcrc_iflg   : out    vl_logic;
        rdusertag_iflg  : out    vl_logic;
        verflut_iflg    : out    vl_logic;
        rdallfault_iflg : out    vl_logic;
        readmfg_iflg    : out    vl_logic;
        vertrim_iflg    : out    vl_logic;
        writecfg_iflg   : out    vl_logic;
        wrrecfg_iflg    : out    vl_logic;
        wrrecfgmask_iflg: out    vl_logic;
        wrallrecfg_iflg : out    vl_logic;
        wrrdvid1_iflg   : out    vl_logic;
        wrrdvid2_iflg   : out    vl_logic;
        wrrdvid3_iflg   : out    vl_logic;
        wrrdvid4_iflg   : out    vl_logic;
        wrrdvid5_iflg   : out    vl_logic;
        wrrdvid6_iflg   : out    vl_logic;
        wrrdvid7_iflg   : out    vl_logic;
        wrrdvid8_iflg   : out    vl_logic;
        writeusertag_iflg: out    vl_logic;
        writemfg_iflg   : out    vl_logic;
        enprog_iflg     : out    vl_logic;
        wri2csa_iflg    : out    vl_logic;
        wrmeasctrl_iflg : out    vl_logic;
        rdmeasresult_iflg: out    vl_logic;
        ldrecfg_pulse   : out    vl_logic;
        wrir_en_i2c_dat : out    vl_logic;
        wr_ir           : out    vl_logic;
        prgmarray       : out    vl_logic;
        noack           : out    vl_logic;
        porsync         : out    vl_logic;
        safestate       : out    vl_logic;
        userlogicrst_pulse: out    vl_logic;
        readtrim_iflg   : out    vl_logic;
        writetrim_iflg  : out    vl_logic;
        rdtrimshdw_iflg : out    vl_logic;
        wrtrimshdw_iflg : out    vl_logic;
        ldtrimshdw_iflg : out    vl_logic;
        rdsoftfault_iflg: out    vl_logic;
        not_verrdall_iflg: out    vl_logic;
        not_rdsoftfault : out    vl_logic;
        m_progcfg_iflg  : out    vl_logic;
        m_progusertag_iflg: out    vl_logic;
        m_progtrim_iflg : out    vl_logic;
        verfault_iflg   : out    vl_logic;
        rdfaulten_iflg  : out    vl_logic;
        tst_north_keeper_iflg: out    vl_logic;
        mc_bus          : in     vl_logic_vector(7 downto 0);
        por             : in     vl_logic;
        reset           : in     vl_logic;
        clk             : in     vl_logic;
        wrir_in         : in     vl_logic;
        refresh_on      : in     vl_logic;
        prgm_mode       : in     vl_logic;
        donebit         : in     vl_logic;
        mfg_mode        : in     vl_logic;
        ld_prgmarray_slaveflgreg: in     vl_logic;
        erase_prgrm_active: in     vl_logic;
        clear_erase_prgrm_flags: in     vl_logic;
        flclr_ep_iflgs  : in     vl_logic;
        ld_rfrsh_sshdw  : in     vl_logic;
        ld_crc_s_latch  : in     vl_logic;
        usertag_enable  : in     vl_logic;
        clear_verrdall_iflg: in     vl_logic;
        clear_rdsoftfault_iflg: in     vl_logic;
        examine_fldonebit: in     vl_logic;
        rst_ldshdw_iflgs: in     vl_logic;
        fsafe           : in     vl_logic
    );
end instruction;
