library verilog;
use verilog.vl_types.all;
entity cfg_logic is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 1;
        DECRYPTION      : integer := 1
    );
    port(
        isc_done        : out    vl_logic;
        lsc_done        : out    vl_logic;
        busy_seldr      : out    vl_logic;
        isc_operational : out    vl_logic;
        jtag_active_smpulse: out    vl_logic;
        jtag_active_smsync: out    vl_logic;
        jtag_active_smsync_jb: out    vl_logic;
        rti2d_smsync    : out    vl_logic;
        rti2d_smpulse   : out    vl_logic;
        jinstr_cap      : out    vl_logic_vector(7 downto 0);
        jconfig_cap     : out    vl_logic_vector(7 downto 0);
        j_com_word4_dat : out    vl_logic_vector(127 downto 0);
        nj_com_word4_dat: out    vl_logic_vector(127 downto 0);
        buf128_int      : out    vl_logic_vector(127 downto 0);
        sector_dat      : out    vl_logic_vector(7 downto 0);
        isc_exec_a      : out    vl_logic;
        isc_exec_b      : out    vl_logic;
        isc_exec_c      : out    vl_logic;
        isc_exec_d      : out    vl_logic;
        isc_exec_e      : out    vl_logic;
        isc_exec_f      : out    vl_logic;
        ref_rst_sync    : out    vl_logic;
        nj_rst_async    : out    vl_logic;
        nj_rst_sync0    : out    vl_logic;
        nj_rst_sync     : out    vl_logic;
        nj_rst_flag     : out    vl_logic;
        nj_rst_ctrl0    : out    vl_logic;
        isc_rst_async   : out    vl_logic;
        isc_rst_sync    : out    vl_logic;
        sf_rst_async    : out    vl_logic;
        sf_rst_sync     : out    vl_logic;
        sed_rst_async   : out    vl_logic;
        sed_rst_sync    : out    vl_logic;
        sed_rst_flag    : out    vl_logic;
        nji2c_rst_async : out    vl_logic;
        njtrx_rst_async : out    vl_logic;
        njtrx_rst_async0: out    vl_logic;
        access_sram     : out    vl_logic;
        access_flash    : out    vl_logic;
        access_tag      : out    vl_logic;
        access_efuse    : out    vl_logic;
        access_sudo     : out    vl_logic;
        access_safe     : out    vl_logic;
        access_mfg      : out    vl_logic;
        access_flash_all: out    vl_logic;
        access_flash_manu: out    vl_logic;
        enter_offline_exec: out    vl_logic;
        enter_offline_eqv: out    vl_logic;
        exit_fl_offline_exec: out    vl_logic;
        exit_normal_exec: out    vl_logic;
        isc_disable_exec: out    vl_logic;
        busy_int        : out    vl_logic;
        fail_int        : out    vl_logic;
        fea_exec_en     : out    vl_logic;
        mfg_margin_en   : out    vl_logic;
        cfg_sed_en      : out    vl_logic;
        sf_prog_sec_eqv : out    vl_logic;
        read_sram_dis   : out    vl_logic;
        write_sram_dis  : out    vl_logic;
        erase_sram_dis  : out    vl_logic;
        read_flfea_dis  : out    vl_logic;
        write_flfea_dis : out    vl_logic;
        erase_flfea_dis : out    vl_logic;
        read_otps_dis   : out    vl_logic;
        write_otps_dis  : out    vl_logic;
        read_flcfg_dis  : out    vl_logic;
        write_flcfg_dis : out    vl_logic;
        erase_flcfg_dis : out    vl_logic;
        read_flufm_dis  : out    vl_logic;
        write_flufm_dis : out    vl_logic;
        erase_flufm_dis : out    vl_logic;
        read_efuse_dis  : out    vl_logic;
        write_efuse_dis : out    vl_logic;
        pwd_mismatch_all: out    vl_logic;
        exec_buf        : out    vl_logic_vector(127 downto 0);
        idcode_err      : out    vl_logic;
        bse_active      : out    vl_logic;
        finish_ppt      : out    vl_logic;
        finish_cdm      : out    vl_logic;
        finish_sdm      : out    vl_logic;
        finish_bke      : out    vl_logic;
        ref_start       : out    vl_logic;
        restart_bse     : out    vl_logic;
        jaccessed_sync  : out    vl_logic;
        burst_start     : out    vl_logic;
        burst_inp       : out    vl_logic;
        jburst_inp      : out    vl_logic;
        dev_sdm_inp     : out    vl_logic;
        restart_bse_en  : out    vl_logic;
        njboot_dat      : out    vl_logic_vector(7 downto 0);
        cib_wkupclk_en  : out    vl_logic;
        cfg_reset_crc16 : out    vl_logic;
        instr_dts       : out    vl_logic;
        start_dts       : out    vl_logic;
        cfg_done_cib    : out    vl_logic;
        gsrn            : out    vl_logic;
        gsrn_sync       : out    vl_logic;
        goe             : out    vl_logic;
        ts_all          : out    vl_logic;
        done_gwe        : out    vl_logic;
        freeze_io       : out    vl_logic;
        freeze_mib      : out    vl_logic;
        pcs_rstn        : out    vl_logic;
        en_pupn         : out    vl_logic;
        stdby_ena       : out    vl_logic;
        dev_stdby_exec  : out    vl_logic;
        dev_sleep_exec  : out    vl_logic;
        dev_wkup_exec   : out    vl_logic;
        dev_sed_exec    : out    vl_logic;
        dev_sdm_qual    : out    vl_logic;
        HFC_EN          : in     vl_logic;
        IDCODE0         : in     vl_logic_vector(31 downto 0);
        CHIPID          : in     vl_logic_vector(7 downto 0);
        por             : in     vl_logic;
        tck             : in     vl_logic;
        smclk           : in     vl_logic;
        hfc_select_pin  : in     vl_logic;
        scanen          : in     vl_logic;
        bg_rdy          : in     vl_logic;
        dts_out         : in     vl_logic_vector(31 downto 0);
        ctrl_nbke       : in     vl_logic;
        ctrl_wkup_tran  : in     vl_logic;
        ctrl_hfc_hd     : in     vl_logic;
        mc1_gsrn_inv    : in     vl_logic;
        mc1_gsrn_sync   : in     vl_logic;
        mc1_user_gsrn   : in     vl_logic;
        mc1_pcs         : in     vl_logic;
        mc1_pupn        : in     vl_logic;
        mc1_en_tsall    : in     vl_logic;
        mc1_tsall_inv   : in     vl_logic;
        mc1_sleep_pupn  : in     vl_logic;
        cib_user_gsr    : in     vl_logic;
        cib_tsall       : in     vl_logic;
        trim_idcode_msb : in     vl_logic_vector(3 downto 0);
        trim_idmsb_en   : in     vl_logic_vector(3 downto 0);
        sed_err         : in     vl_logic;
        sed_busy        : in     vl_logic;
        sed_active      : in     vl_logic;
        sed_boot        : in     vl_logic;
        programn_tog    : in     vl_logic;
        gsrn_pin_sync   : in     vl_logic;
        boot_setup      : in     vl_logic_vector(5 downto 0);
        wbc_active      : in     vl_logic;
        ref_states      : in     vl_logic_vector(6 downto 0);
        ref_dones       : in     vl_logic_vector(5 downto 0);
        ref_ppt         : in     vl_logic;
        ref_cdm         : in     vl_logic;
        exit_accessed   : in     vl_logic;
        initn_tmr       : in     vl_logic;
        wkup_done       : in     vl_logic;
        wkup_done_rise  : in     vl_logic;
        gsrn_tmr        : in     vl_logic;
        gwe_tmr         : in     vl_logic;
        goe_tmr         : in     vl_logic;
        fio_tmr         : in     vl_logic;
        fmib_tmr        : in     vl_logic;
        wkup_aux_pulse  : in     vl_logic;
        sleep_mode_flag : in     vl_logic;
        wkup_done_cib   : in     vl_logic;
        lsc_sdm         : in     vl_logic;
        bsmode1         : in     vl_logic;
        tsall_ctrl      : in     vl_logic;
        isc_enabled     : in     vl_logic;
        isc_disable_completing: in     vl_logic;
        jset_isc_done_i : in     vl_logic;
        jrst_isc_done_i : in     vl_logic;
        jtag_active     : in     vl_logic;
        rti2d           : in     vl_logic;
        seldr_ss        : in     vl_logic;
        capdr_ss_r      : in     vl_logic;
        jaccess_sram    : in     vl_logic;
        jaccess_flash   : in     vl_logic;
        jaccess_fl_norm : in     vl_logic;
        jaccess_fl_sudo : in     vl_logic;
        jaccess_fl_safe : in     vl_logic;
        jaccess_efuse   : in     vl_logic;
        jaccess_ef_norm : in     vl_logic;
        jaccess_ef_sudo : in     vl_logic;
        jaccess_ef_safe : in     vl_logic;
        jaccess_tag     : in     vl_logic;
        jaccess_flash_all: in     vl_logic;
        jenable_offl    : in     vl_logic;
        jconfig_dat     : in     vl_logic_vector(3 downto 0);
        jsector_dat     : in     vl_logic_vector(7 downto 0);
        jbuf128_dat     : in     vl_logic_vector(127 downto 0);
        j_enable_qual   : in     vl_logic;
        j_enable_x_qual : in     vl_logic;
        j_disable_qual  : in     vl_logic;
        jexit_fl_offline: in     vl_logic;
        jexit_normal    : in     vl_logic;
        mfg_en          : in     vl_logic;
        mfg_margin      : in     vl_logic;
        mfg_bkgrndft_en : in     vl_logic;
        jburst_en       : in     vl_logic;
        isc_nj_enabled  : in     vl_logic;
        isc_nj_disable_completing: in     vl_logic;
        njset_isc_done_c: in     vl_logic;
        njrst_isc_done_c: in     vl_logic;
        njtag_active    : in     vl_logic;
        njtag_active_nsed: in     vl_logic;
        njaccess_sram   : in     vl_logic;
        njaccess_flash  : in     vl_logic;
        njaccess_fl_norm: in     vl_logic;
        njaccess_fl_sudo: in     vl_logic;
        njaccess_fl_safe: in     vl_logic;
        njaccess_efuse  : in     vl_logic;
        njaccess_ef_norm: in     vl_logic;
        njaccess_ef_sudo: in     vl_logic;
        njaccess_ef_safe: in     vl_logic;
        njaccess_tag    : in     vl_logic;
        njaccess_flash_all: in     vl_logic;
        njenable_offl   : in     vl_logic;
        nj_exec_a       : in     vl_logic;
        nj_exec_b       : in     vl_logic;
        nj_exec_c       : in     vl_logic;
        nj_exec_d       : in     vl_logic;
        nj_exec_e       : in     vl_logic;
        nj_exec_f       : in     vl_logic;
        njconfig_dat    : in     vl_logic_vector(3 downto 0);
        njsector_dat    : in     vl_logic_vector(7 downto 0);
        njbuf128_dat    : in     vl_logic_vector(127 downto 0);
        nj_enable_qual  : in     vl_logic;
        nj_enable_x_qual: in     vl_logic;
        nj_disable_qual : in     vl_logic;
        njexit_fl_offline: in     vl_logic;
        njexit_normal   : in     vl_logic;
        njburst_inp     : in     vl_logic;
        njbse_init      : in     vl_logic;
        njbse_txcmd     : in     vl_logic;
        njbse_preamble  : in     vl_logic;
        njbse_rxcmd     : in     vl_logic;
        njbse_rxdec     : in     vl_logic;
        njbse_bypass    : in     vl_logic;
        njbse_fthrough  : in     vl_logic;
        finish_bse      : in     vl_logic;
        njbse_err_bus   : in     vl_logic_vector(3 downto 0);
        preamble_std    : in     vl_logic;
        preamble_enc    : in     vl_logic;
        mstr_busy_bse   : in     vl_logic;
        sd_sram_otp     : in     vl_logic;
        sd_fea_otp      : in     vl_logic;
        sd_cfg_otp      : in     vl_logic;
        sd_ufm_otp      : in     vl_logic;
        sd_key_lock     : in     vl_logic;
        sd_dec_only     : in     vl_logic;
        sd_pwd_mismatch : in     vl_logic;
        sd_assp_en      : in     vl_logic;
        sd_pwd_en       : in     vl_logic;
        sd_pwd_all      : in     vl_logic;
        sd_red_en       : in     vl_logic;
        sd_red_plc      : in     vl_logic;
        sd_red_ebr      : in     vl_logic;
        ctrl0           : in     vl_logic_vector(31 downto 0);
        cidcode         : in     vl_logic_vector(31 downto 0);
        uidcode         : in     vl_logic_vector(63 downto 0);
        comp_dic        : in     vl_logic_vector(63 downto 0);
        cfg_reg_dat     : in     vl_logic_vector(127 downto 0);
        cfg_crc         : in     vl_logic_vector(15 downto 0);
        mt_freq_cnt     : in     vl_logic_vector(15 downto 0);
        id_err          : in     vl_logic;
        njs_invalid_err : in     vl_logic;
        sram_sec_prog   : in     vl_logic;
        sram_sec_read   : in     vl_logic;
        sram_done       : in     vl_logic;
        sram_ues        : in     vl_logic_vector(31 downto 0);
        sf_exec_buf     : in     vl_logic_vector(127 downto 0);
        busy_sram       : in     vl_logic;
        fail_sram       : in     vl_logic;
        sf_finish_bke   : in     vl_logic;
        flash_sec_prog  : in     vl_logic;
        flash_sec_read  : in     vl_logic;
        flash_secplus   : in     vl_logic;
        flash_done      : in     vl_logic;
        flash_ues       : in     vl_logic_vector(31 downto 0);
        fl_exec_buf     : in     vl_logic_vector(127 downto 0);
        fl_modal_state  : in     vl_logic_vector(31 downto 0);
        fl_pg_count     : in     vl_logic_vector(9 downto 0);
        fl_er_count     : in     vl_logic_vector(11 downto 0);
        row             : in     vl_logic_vector(14 downto 6);
        busy_flash      : in     vl_logic;
        fail_flash      : in     vl_logic;
        fl_busy_ppt     : in     vl_logic;
        fl_busy_cdm     : in     vl_logic;
        fl_busy_sdm     : in     vl_logic;
        fl_finish_ppt   : in     vl_logic;
        fl_finish_cdm   : in     vl_logic;
        fl_finish_sdm   : in     vl_logic;
        ef_exec_buf     : in     vl_logic_vector(127 downto 0);
        busy_efuse      : in     vl_logic;
        fail_efuse      : in     vl_logic;
        ef_busy_ppt     : in     vl_logic;
        ef_busy_cdm     : in     vl_logic;
        ef_finish_ppt   : in     vl_logic;
        ef_finish_cdm   : in     vl_logic;
        busy_bse        : in     vl_logic;
        busy_wkup       : in     vl_logic;
        fail_bse        : in     vl_logic;
        lsc_refresh_iq  : in     vl_logic;
        lsc_refresh_cq  : in     vl_logic;
        lsc_jump_cq     : in     vl_logic;
        lsc_chip_select_cq: in     vl_logic;
        verify_id_qual  : in     vl_logic;
        read_temp_qual  : in     vl_logic;
        idcode_pub_iq   : in     vl_logic;
        idcode_prv_iq   : in     vl_logic;
        uidcode_pub_iq  : in     vl_logic;
        usercode_iq     : in     vl_logic;
        read_temp_iq    : in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic;
        lsc_read_status_mq: in     vl_logic;
        lsc_read_mfg_status_mq: in     vl_logic;
        mfg_mdata_mq    : in     vl_logic;
        idcode_pub_cq   : in     vl_logic;
        idcode_prv_cq   : in     vl_logic;
        uidcode_pub_cq  : in     vl_logic;
        usercode_cq     : in     vl_logic;
        read_temp_cq    : in     vl_logic;
        lsc_read_status_cq: in     vl_logic;
        lsc_check_busy_cq: in     vl_logic;
        lsc_bitstream_burst_qual: in     vl_logic;
        lsc_read_ctrl0_qual: in     vl_logic;
        lsc_read_crc_qual: in     vl_logic;
        lsc_read_comp_dic_qual: in     vl_logic;
        lsc_reset_crc_qual: in     vl_logic;
        sf_prog_std_all : in     vl_logic;
        sf_prog_enc_all : in     vl_logic;
        lsc_device_ctrl_qual: in     vl_logic;
        fl_erase_qual   : in     vl_logic;
        fl_erase_tag_qual: in     vl_logic;
        cmd_read_exec_buf: in     vl_logic;
        cmd_prog_cfg_reg: in     vl_logic;
        cmd_read_cfg_reg: in     vl_logic;
        lsc_read_i2c_qual: in     vl_logic;
        cfg_i2c_dout    : in     vl_logic_vector(7 downto 0)
    );
end cfg_logic;
