library verilog;
use verilog.vl_types.all;
entity ser_aux_top is
    port(
        atsten          : out    vl_logic;
        bitclk_from_nd_eno: out    vl_logic;
        bs4refck        : out    vl_logic;
        bus8bit_selo    : out    vl_logic;
        cdr_lol_setvcc  : out    vl_logic_vector(1 downto 0);
        ck3g4txn        : out    vl_logic;
        ck3g4txn2nd     : out    vl_logic;
        ck3g4txp        : out    vl_logic;
        ck3g4txp2nd     : out    vl_logic;
        dco_calib_time_selvcc: out    vl_logic_vector(1 downto 0);
        iref_50uconst_ch: out    vl_logic_vector(3 downto 0);
        iref_50urpoly_ch: out    vl_logic_vector(3 downto 0);
        isetloso        : out    vl_logic_vector(7 downto 0);
        lol_div_vcc     : out    vl_logic_vector(1 downto 0);
        macropdbvcc     : out    vl_logic;
        pd_iseto        : out    vl_logic_vector(1 downto 0);
        plol            : out    vl_logic;
        plol_sts        : out    vl_logic;
        plol_stsb       : out    vl_logic;
        refck2core      : out    vl_logic;
        refck25xo       : out    vl_logic;
        refck_modeo     : out    vl_logic_vector(1 downto 0);
        refck2ndp       : out    vl_logic;
        refck2ndn       : out    vl_logic;
        reg2fpga_out    : out    vl_logic;
        req_iseto       : out    vl_logic_vector(2 downto 0);
        reset_vcc       : out    vl_logic;
        reseto          : out    vl_logic;
        rx_bs_modeo     : out    vl_logic;
        rx_refck_local  : out    vl_logic;
        seticonst_cho   : out    vl_logic_vector(1 downto 0);
        setirpoly_cho   : out    vl_logic_vector(1 downto 0);
        sync            : out    vl_logic;
        sync_local_eno  : out    vl_logic;
        sync_nd_eno     : out    vl_logic;
        sync_pulse2ndp  : out    vl_logic;
        sync_pulse2ndn  : out    vl_logic;
        tck_full        : out    vl_logic;
        tielow_aux      : out    vl_logic;
        tx_bs_modeo     : out    vl_logic;
        zero            : out    vl_logic_vector(7 downto 0);
        atstn           : inout  vl_logic;
        atstp           : inout  vl_logic;
        iref_50uconst   : inout  vl_logic_vector(1 downto 0);
        iref_50urpoly   : inout  vl_logic_vector(1 downto 0);
        vcc             : inout  vl_logic;
        vcca            : inout  vl_logic;
        vcca25          : inout  vl_logic;
        vss             : inout  vl_logic;
        vssa            : inout  vl_logic;
        aux_spare_inb   : in     vl_logic_vector(7 downto 0);
        bitclk_from_nd_en: in     vl_logic;
        bitclk_local_en : in     vl_logic;
        bitclk_nd_en    : in     vl_logic;
        bus8bit_sel     : in     vl_logic;
        cdr_lol_set     : in     vl_logic_vector(1 downto 0);
        ck_core_tx      : in     vl_logic;
        cmusetbiasi     : in     vl_logic_vector(1 downto 0);
        dco_calib_time_sel: in     vl_logic_vector(1 downto 0);
        ib_pwdnb        : in     vl_logic;
        isetlos         : in     vl_logic_vector(7 downto 0);
        lol_div         : in     vl_logic_vector(1 downto 0);
        macropdb        : in     vl_logic;
        macrorst        : in     vl_logic;
        pd_iset         : in     vl_logic_vector(1 downto 0);
        pll_lol_set     : in     vl_logic_vector(1 downto 0);
        pwr_on_rst      : in     vl_logic;
        refck25x        : in     vl_logic;
        refck_dcbias_en : in     vl_logic;
        refck_from_nd   : in     vl_logic;
        refck_from_nd_sel: in     vl_logic_vector(1 downto 0);
        refck_mode      : in     vl_logic_vector(1 downto 0);
        refck_out_sel   : in     vl_logic_vector(1 downto 0);
        refck_pwdnb     : in     vl_logic;
        refck_rterm     : in     vl_logic;
        refck_to_nd_en  : in     vl_logic;
        refclkn         : in     vl_logic;
        refclkp         : in     vl_logic;
        reg2fpga_ctrl   : in     vl_logic;
        req_iset        : in     vl_logic_vector(2 downto 0);
        rg_en           : in     vl_logic;
        rg_set          : in     vl_logic_vector(1 downto 0);
        rx_bs_mode      : in     vl_logic;
        rx_hstest1      : in     vl_logic_vector(1 downto 0);
        rx_lstest1      : in     vl_logic_vector(1 downto 0);
        rx_lstest2      : in     vl_logic_vector(1 downto 0);
        rx_lstest3      : in     vl_logic_vector(1 downto 0);
        ser_mem         : in     vl_logic_vector(41 downto 8);
        seticonst_aux   : in     vl_logic_vector(1 downto 0);
        seticonst_ch    : in     vl_logic_vector(1 downto 0);
        setirpoly_aux   : in     vl_logic_vector(1 downto 0);
        setirpoly_ch    : in     vl_logic_vector(1 downto 0);
        setpllrc        : in     vl_logic_vector(5 downto 0);
        sync_local_en   : in     vl_logic;
        sync_nd_en      : in     vl_logic;
        sync_pulse      : in     vl_logic;
        trst            : in     vl_logic;
        tst_en          : in     vl_logic;
        tst_sel         : in     vl_logic_vector(3 downto 0);
        tx_bs_mode      : in     vl_logic;
        tx_refck_sel    : in     vl_logic;
        tx_vco_ck_div   : in     vl_logic_vector(2 downto 0);
        txpll_pwdnb     : in     vl_logic
    );
end ser_aux_top;
