library verilog;
use verilog.vl_types.all;
entity cfg_register is
    generic(
        FLASH_MEM       : integer := 1;
        EFUSE_MEM       : integer := 1;
        DECRYPTION      : integer := 1
    );
    port(
        fsd_persistn_progn: out    vl_logic;
        fsd_persist_initn: out    vl_logic;
        fsd_persist_done: out    vl_logic;
        fsd_persistn_jtag: out    vl_logic;
        fsd_persistn_sspi: out    vl_logic;
        fsd_persistn_i2c: out    vl_logic;
        fsd_persist_mspi: out    vl_logic;
        fsd_boot_sel    : out    vl_logic_vector(1 downto 0);
        fsd_gold_addr   : out    vl_logic_vector(15 downto 0);
        sd_i2c_addr     : out    vl_logic_vector(7 downto 0);
        sd_key_lock     : out    vl_logic;
        sd_dec_only     : out    vl_logic;
        sd_pwd_en       : out    vl_logic;
        sd_pwd_all      : out    vl_logic;
        sd_assp_en      : out    vl_logic;
        sd_sram_otp     : out    vl_logic;
        sd_fea_otp      : out    vl_logic;
        sd_cfg_otp      : out    vl_logic;
        sd_ufm_otp      : out    vl_logic;
        sd_pwd_mismatch : out    vl_logic;
        sd_red_en       : out    vl_logic;
        sd_red_plc      : out    vl_logic;
        sd_red_ebr      : out    vl_logic;
        sd_trim         : out    vl_logic_vector(127 downto 0);
        ctrl0           : out    vl_logic_vector(31 downto 0);
        cidcode         : out    vl_logic_vector(31 downto 0);
        uidcode         : out    vl_logic_vector(63 downto 0);
        comp_dic        : out    vl_logic_vector(63 downto 0);
        sd_key_last     : out    vl_logic_vector(127 downto 0);
        mt_freq_cnt     : out    vl_logic_vector(15 downto 0);
        cfg_reg_dat     : out    vl_logic_vector(127 downto 0);
        id_err          : out    vl_logic;
        njs_invalid_err : out    vl_logic;
        buf128_dat      : out    vl_logic_vector(127 downto 0);
        cfg_i2c_dat     : out    vl_logic_vector(15 downto 0);
        cfg_ctrl0_upd   : out    vl_logic;
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        nj_rst_flag     : in     vl_logic;
        scanen          : in     vl_logic;
        CTRL0_DEFAULT   : in     vl_logic_vector(31 downto 0);
        ASSP_EN         : in     vl_logic;
        ENC_ONLY_EN     : in     vl_logic;
        p_slave         : in     vl_logic;
        bg_cmp_out      : in     vl_logic;
        proc_ring_osc   : in     vl_logic;
        mfg_freq_sel    : in     vl_logic;
        mfg_bkgrndft_en : in     vl_logic;
        buf128_int      : in     vl_logic_vector(127 downto 0);
        sector_dat      : in     vl_logic_vector(7 downto 0);
        nj_exec_b       : in     vl_logic;
        isc_exec_e      : in     vl_logic;
        idcode_err      : in     vl_logic;
        bse_active      : in     vl_logic;
        mfg_en          : in     vl_logic;
        access_sudo     : in     vl_logic;
        access_safe     : in     vl_logic;
        rti_r           : in     vl_logic;
        upir_ss_r       : in     vl_logic;
        exit1dr_ss_r    : in     vl_logic;
        ref_start       : in     vl_logic;
        nj_rst_ctrl0    : in     vl_logic;
        rst_ctrl0_onfail: in     vl_logic;
        bse_err_rst     : in     vl_logic;
        access_flash_manu: in     vl_logic;
        fl_load_trim    : in     vl_logic;
        fl_load_pes     : in     vl_logic;
        fl_load_mes     : in     vl_logic;
        fl_load_key     : in     vl_logic;
        fl_load_pwd     : in     vl_logic;
        fl_load_fea     : in     vl_logic;
        fl_load_feabits : in     vl_logic;
        fl_load_otps    : in     vl_logic;
        fl_erase_trim   : in     vl_logic;
        fl_erase_fea    : in     vl_logic;
        ef_load_trim    : in     vl_logic;
        ef_load_pes     : in     vl_logic;
        ef_load_mes     : in     vl_logic;
        ef_load_key     : in     vl_logic;
        ef_load_pwd     : in     vl_logic;
        ef_load_fea     : in     vl_logic;
        ef_load_feabits : in     vl_logic;
        ef_load_otps    : in     vl_logic;
        verify_id_qual  : in     vl_logic;
        lsc_prog_ctrl0_qual: in     vl_logic;
        lsc_write_comp_dic_qual: in     vl_logic;
        lsc_shift_password_qual: in     vl_logic;
        isc_prog_done_qual: in     vl_logic;
        isc_prog_sec_qual: in     vl_logic;
        isc_prog_secplus_qual: in     vl_logic;
        lsc_prog_password_qual: in     vl_logic;
        lsc_prog_cipher_key_qual: in     vl_logic;
        lsc_prog_feature_qual: in     vl_logic;
        lsc_prog_feabits_qual: in     vl_logic;
        lsc_prog_otps_qual: in     vl_logic;
        lsc_prog_trim_qual: in     vl_logic;
        lsc_prog_pes_qual: in     vl_logic;
        lsc_prog_mes_qual: in     vl_logic;
        lsc_read_password_qual: in     vl_logic;
        lsc_read_cipher_key_qual: in     vl_logic;
        lsc_read_feature_qual: in     vl_logic;
        lsc_read_feabits_qual: in     vl_logic;
        lsc_read_otps_qual: in     vl_logic;
        lsc_read_trim_qual: in     vl_logic;
        lsc_read_pes_qual: in     vl_logic;
        lsc_read_mes_qual: in     vl_logic;
        fl_write_addr_qual: in     vl_logic;
        mfg_mdata_qual  : in     vl_logic;
        mfg_mtrim_qual  : in     vl_logic;
        sed_prog_ctrl0_qual: in     vl_logic;
        sed_write_comp_dic_qual: in     vl_logic;
        isc_disable_exec: in     vl_logic;
        exec_buf        : in     vl_logic_vector(127 downto 0);
        njs_invalid_c   : in     vl_logic
    );
end cfg_register;
