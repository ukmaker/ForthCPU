library verilog;
use verilog.vl_types.all;
entity datap_unit is
    generic(
        DECRYPTION      : integer := 1
    );
    port(
        njtag_run       : out    vl_logic;
        nj_dat_ren      : out    vl_logic;
        nj_dat_wen      : out    vl_logic;
        njtag_din       : out    vl_logic_vector(7 downto 0);
        decompress_njtag_en: out    vl_logic;
        dec_load        : out    vl_logic;
        rfifo_re        : out    vl_logic;
        wfifo_we        : out    vl_logic;
        wfifo_din       : out    vl_logic_vector(7 downto 0);
        decompress_1byte: out    vl_logic;
        decompress_8byte: out    vl_logic;
        decompress_out  : out    vl_logic_vector(63 downto 0);
        decrypt_burst   : out    vl_logic;
        decrypt_out     : out    vl_logic_vector(7 downto 0);
        dp_dsr_8byte_cmp: out    vl_logic;
        dp_dsr_1byte_cmp: out    vl_logic;
        dp_dsr_1byte_enc: out    vl_logic;
        cfg_crc         : out    vl_logic_vector(15 downto 0);
        njm_crc_err     : out    vl_logic;
        sdm_run         : out    vl_logic;
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        isc_rst_sync    : in     vl_logic;
        sed_en_adv      : in     vl_logic;
        sed_active      : in     vl_logic;
        njtag_slv_en    : in     vl_logic;
        njfsm_hold      : in     vl_logic;
        jtag_active_smsync: in     vl_logic;
        ShiftDR         : in     vl_logic;
        isc_data_shift_iqual: in     vl_logic;
        lsc_prog_incr_rti_iqual: in     vl_logic;
        lsc_prog_incr_enc_iqual: in     vl_logic;
        lsc_prog_incr_cne_iqual: in     vl_logic;
        lsc_prog_incr_cmp_iqual: in     vl_logic;
        lsc_bitstream_burst_iq: in     vl_logic;
        njtag_active    : in     vl_logic;
        njtag_cmd       : in     vl_logic;
        njtag_infa      : in     vl_logic;
        njshf_dat0      : in     vl_logic;
        njshf_dat       : in     vl_logic;
        njshf_crc       : in     vl_logic;
        njshf_dum       : in     vl_logic;
        njbse_rxcmd     : in     vl_logic;
        njbse_rxdec     : in     vl_logic;
        isc_data_shift_cqual: in     vl_logic;
        lsc_prog_incr_rti_cqual: in     vl_logic;
        lsc_prog_incr_enc_cqual: in     vl_logic;
        lsc_prog_incr_cne_cqual: in     vl_logic;
        lsc_prog_incr_cmp_cqual: in     vl_logic;
        nj_cmd_read_com : in     vl_logic;
        nj_cmd_read_dsr : in     vl_logic;
        nj_cmd_prog_com : in     vl_logic;
        j_ins_prog_com  : in     vl_logic;
        jburst_inp      : in     vl_logic;
        dev_sdm_inp     : in     vl_logic;
        cfg_reset_crc16 : in     vl_logic;
        nj_check_crc    : in     vl_logic;
        decom_last_mask : in     vl_logic;
        dum_dat         : in     vl_logic_vector(7 downto 0);
        jbuf8_rdy       : in     vl_logic;
        jbuf8_dat       : in     vl_logic_vector(7 downto 0);
        njcom_out       : in     vl_logic_vector(7 downto 0);
        dsr_out         : in     vl_logic_vector(7 downto 0);
        wfifo_full      : in     vl_logic;
        rfifo_empty     : in     vl_logic;
        rfifo_out       : in     vl_logic_vector(7 downto 0);
        sd_key_last     : in     vl_logic_vector(127 downto 0);
        comp_dic        : in     vl_logic_vector(63 downto 0);
        lsc_sdm         : in     vl_logic;
        dnld_dat        : in     vl_logic_vector(7 downto 0);
        dnld_dat_en     : in     vl_logic
    );
end datap_unit;
