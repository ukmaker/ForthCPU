library verilog;
use verilog.vl_types.all;
entity cfg_bse is
    generic(
        st_idle         : integer := 0;
        st_init         : integer := 1;
        st_rstsst       : integer := 3;
        st_postrst      : integer := 7;
        st_setsst       : integer := 5;
        st_postsst      : integer := 14;
        st_setmp        : integer := 9;
        st_txcmd        : integer := 13;
        st_preamble     : integer := 15;
        st_rxcmd        : integer := 12;
        st_rxdec        : integer := 6;
        st_bypass       : integer := 11;
        st_fthrough     : integer := 10;
        st_error        : integer := 2;
        st_finish       : integer := 4;
        st_abort        : integer := 8;
        setup_idle      : integer := 0;
        setup_init      : integer := 1;
        setup_mcpu      : integer := 3;
        setup_mcmd      : integer := 5;
        setup_mop1      : integer := 7;
        setup_mop2      : integer := 6;
        setup_mop3      : integer := 4;
        setup_done      : integer := 2
    );
    port(
        njbse_init      : out    vl_logic;
        njbse_sstcmd    : out    vl_logic;
        njbse_txcmd     : out    vl_logic;
        njbse_preamble  : out    vl_logic;
        njbse_rxcmd     : out    vl_logic;
        njbse_rxdec     : out    vl_logic;
        njbse_rxall     : out    vl_logic;
        njbse_bypass    : out    vl_logic;
        njbse_fthrough  : out    vl_logic;
        cfg_mstr_start  : out    vl_logic;
        cfg_mstr_stop   : out    vl_logic;
        tx_setmcpu      : out    vl_logic;
        tx_command      : out    vl_logic;
        tx_operand      : out    vl_logic;
        cfg_mtx_dat     : out    vl_logic_vector(7 downto 0);
        cfg_mcsn_dat    : out    vl_logic_vector(7 downto 0);
        busy_bse        : out    vl_logic;
        fail_bse        : out    vl_logic;
        finish_bse      : out    vl_logic;
        bse_err_rst     : out    vl_logic;
        njbse_err_bus   : out    vl_logic_vector(3 downto 0);
        mstr_busy_bse   : out    vl_logic;
        last_addr_cib   : out    vl_logic_vector(15 downto 0);
        nj_rst_async    : in     vl_logic;
        nj_rst_sync0    : in     vl_logic;
        nj_rst_flag     : in     vl_logic;
        smclk           : in     vl_logic;
        ctrl_mspim_sel  : in     vl_logic;
        ctrl_pdone_ovld : in     vl_logic_vector(1 downto 0);
        cib_mspim_addr  : in     vl_logic_vector(15 downto 0);
        cib_mcsn_sel    : in     vl_logic;
        mc1_mspi_sed_addr: in     vl_logic_vector(15 downto 0);
        mc1_source_sel  : in     vl_logic;
        mc1_mspi_addr   : in     vl_logic_vector(15 downto 0);
        p_slave         : in     vl_logic;
        p_mspi0         : in     vl_logic;
        p_mspim         : in     vl_logic;
        p_mp8           : in     vl_logic;
        p_mp16          : in     vl_logic;
        p_mspi_slow     : in     vl_logic;
        p_mspi_fast     : in     vl_logic;
        p_mspi_dual     : in     vl_logic;
        p_mspi_quad     : in     vl_logic;
        p_mp8_quad      : in     vl_logic;
        p_mp16_quad     : in     vl_logic;
        p_mspi_all      : in     vl_logic;
        p_sst           : in     vl_logic;
        p_end_bpft      : in     vl_logic;
        done_rise1      : in     vl_logic;
        start_bse0      : in     vl_logic;
        start_bse1      : in     vl_logic;
        start_bse2      : in     vl_logic;
        int_prm_nrdy    : in     vl_logic;
        ref_boot1       : in     vl_logic;
        cfg_mstr_busy   : in     vl_logic;
        njm_tr_next     : in     vl_logic;
        njm_tr_done     : in     vl_logic;
        njm_mcpu_done   : in     vl_logic;
        preamble_std    : in     vl_logic;
        preamble_enc    : in     vl_logic;
        preamble_err    : in     vl_logic;
        lsc_jump_cq     : in     vl_logic;
        lsc_chip_select_cq: in     vl_logic;
        jump_exec       : in     vl_logic;
        chip_select_exec: in     vl_logic;
        flow_through_exec: in     vl_logic;
        bypass_exec     : in     vl_logic;
        bse_end_cqual   : in     vl_logic;
        bse_prog_incr_cqual: in     vl_logic;
        njm_invalid_c   : in     vl_logic;
        njr_invalid_c   : in     vl_logic;
        sed_invalid_c   : in     vl_logic;
        nj_jump_param   : in     vl_logic_vector(31 downto 0);
        nj_csel_param   : in     vl_logic_vector(7 downto 0);
        nj_exec_b       : in     vl_logic;
        njm_crc_err     : in     vl_logic;
        id_err          : in     vl_logic;
        burst_start     : in     vl_logic;
        burst_inp       : in     vl_logic;
        sd_dec_only     : in     vl_logic;
        restart_bse     : in     vl_logic;
        ref_start       : in     vl_logic;
        sed_en_adv      : in     vl_logic;
        sed_start_bse   : in     vl_logic;
        lsc_sdm         : in     vl_logic;
        sdm_start_bse   : in     vl_logic;
        sdm_bse_eof     : in     vl_logic;
        preamble_std_sdm: in     vl_logic;
        preamble_enc_sdm: in     vl_logic;
        preamble_err_sdm: in     vl_logic;
        sf_asr_out      : in     vl_logic
    );
end cfg_bse;
