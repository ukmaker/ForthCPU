library verilog;
use verilog.vl_types.all;
entity invx8v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end invx8v1s;
