library verilog;
use verilog.vl_types.all;
entity pcs_or2_2 is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        X               : out    vl_logic
    );
end pcs_or2_2;
