library verilog;
use verilog.vl_types.all;
entity cfg_driver is
    port(
        dsr_clk         : out    vl_logic;
        dsr_din         : out    vl_logic_vector(63 downto 0);
        dsr_shift       : out    vl_logic_vector(1 downto 0);
        dsr_rst_n       : out    vl_logic;
        dsr_cap         : out    vl_logic;
        dsr_upd_lat     : out    vl_logic;
        dsr_cnt_en      : out    vl_logic;
        sram_asr_clk    : out    vl_logic;
        sram_asr_in     : out    vl_logic;
        sram_asr_rst    : out    vl_logic;
        sram_asr_en_incr: out    vl_logic;
        sram_asr_shift_1st: out    vl_logic;
        sram_asr_shift_2nd: out    vl_logic;
        sram_asr_shift_3rd: out    vl_logic;
        sram_wl_str     : out    vl_logic;
        sram_data_wr    : out    vl_logic;
        es_o            : out    vl_logic_vector(35 downto 0);
        pcs_o           : out    vl_logic_vector(27 downto 0);
        sed_adv_shf     : out    vl_logic;
        sed_adv_mask    : out    vl_logic_vector(7 downto 0);
        tdrclk          : in     vl_logic;
        dsr_out         : in     vl_logic_vector(7 downto 0);
        ShiftDR         : in     vl_logic;
        ins_dsr_1bit    : in     vl_logic;
        ins_dsr_1byte   : in     vl_logic;
        tdi_dsr_1bit    : in     vl_logic;
        tdi_dsr_1byte   : in     vl_logic_vector(7 downto 0);
        jsel_sram_asr   : in     vl_logic;
        cmd_dsr_1byte   : in     vl_logic;
        nj_dsr_shf      : in     vl_logic;
        nj_dsr_data     : in     vl_logic_vector(7 downto 0);
        decompress_1byte: in     vl_logic;
        decompress_8byte: in     vl_logic;
        decompress_out  : in     vl_logic_vector(63 downto 0);
        decrypt_burst   : in     vl_logic;
        decrypt_out     : in     vl_logic_vector(7 downto 0);
        dp_dsr_8byte_cmp: in     vl_logic;
        dp_dsr_1byte_cmp: in     vl_logic;
        dp_dsr_1byte_enc: in     vl_logic;
        sed_dsr_loop_en : in     vl_logic;
        sed_dsr_1byte   : in     vl_logic;
        tdi_sram_asr    : in     vl_logic;
        sf_dsr_rst      : in     vl_logic;
        sf_dsr_cap      : in     vl_logic;
        sf_dsr_upd_lat  : in     vl_logic;
        sf_asr_in       : in     vl_logic;
        sf_asr_rst      : in     vl_logic;
        sf_asr_en_incr  : in     vl_logic;
        sf_asr_shift_1st: in     vl_logic;
        sf_asr_shift_2nd: in     vl_logic;
        sf_asr_shift_3rd: in     vl_logic;
        sf_wl_str       : in     vl_logic;
        sf_data_wr      : in     vl_logic;
        sf_es_o         : in     vl_logic_vector(35 downto 0);
        sf_pcs_o        : in     vl_logic_vector(27 downto 0);
        ppt_dat         : in     vl_logic_vector(7 downto 0);
        ppt_dsr_shf8_en : in     vl_logic;
        ppt_dsr_shf     : in     vl_logic
    );
end cfg_driver;
