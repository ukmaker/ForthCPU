library verilog;
use verilog.vl_types.all;
entity jtag_register is
    port(
        instruction     : out    vl_logic_vector(7 downto 0);
        ir_sr           : out    vl_logic_vector(7 downto 0);
        jconfig_dat     : out    vl_logic_vector(3 downto 0);
        jsector_dat     : out    vl_logic_vector(7 downto 0);
        jbuf8_rdy       : out    vl_logic;
        jbuf8_dat       : out    vl_logic_vector(7 downto 0);
        jbuf128_dat     : out    vl_logic_vector(127 downto 0);
        mfg_dat         : out    vl_logic_vector(119 downto 0);
        mfg_en          : out    vl_logic;
        tdo_out         : out    vl_logic;
        tdo_oe_out      : out    vl_logic;
        tdi_dsr_1bit    : out    vl_logic;
        tdi_dsr_1byte   : out    vl_logic_vector(7 downto 0);
        tdi_sram_asr    : out    vl_logic;
        tdi_bscan       : out    vl_logic;
        tdi_iscan       : out    vl_logic;
        jpspi_ctrl      : out    vl_logic_vector(15 downto 0);
        por             : in     vl_logic;
        tck             : in     vl_logic;
        tdi             : in     vl_logic;
        tms             : in     vl_logic;
        tlreset         : in     vl_logic;
        selir_ss        : in     vl_logic;
        capir_ss        : in     vl_logic;
        exit1ir_ss      : in     vl_logic;
        exit2ir_ss      : in     vl_logic;
        upir_ss         : in     vl_logic;
        capdr_ss        : in     vl_logic;
        updr_ss         : in     vl_logic;
        ShiftIR         : in     vl_logic;
        ShiftDR         : in     vl_logic;
        jtag_ir_access  : in     vl_logic;
        jsel_byp        : in     vl_logic;
        jsel_cfg        : in     vl_logic;
        jsel_sec        : in     vl_logic;
        jsel_com        : in     vl_logic;
        jsel_com_lsbf   : in     vl_logic;
        jsel_com_msbf   : in     vl_logic;
        jcap_com_word4  : in     vl_logic;
        jshf_com_byte1  : in     vl_logic;
        jshf_com_byte1_msbf: in     vl_logic;
        jshf_com_byte2  : in     vl_logic;
        jshf_com_byte4  : in     vl_logic;
        jshf_com_byte8  : in     vl_logic;
        jshf_com_byte9_msbf: in     vl_logic;
        jshf_com_word4  : in     vl_logic;
        jshf_com_word4_msbf: in     vl_logic;
        jbuf8_s01       : in     vl_logic;
        jbuf8_p08       : in     vl_logic;
        jbuf8_rst       : in     vl_logic;
        jsel_busy       : in     vl_logic;
        jsel_er1        : in     vl_logic;
        jsel_er2        : in     vl_logic;
        jsel_bsr        : in     vl_logic;
        jsel_sram_asr   : in     vl_logic;
        jsel_dsr        : in     vl_logic;
        jsel_mfg        : in     vl_logic;
        jsel_iscan      : in     vl_logic;
        jsel_extspi_i   : in     vl_logic;
        jsel_extspi     : in     vl_logic;
        lsc_iscan_m     : in     vl_logic_vector(7 downto 0);
        j_enable_qual   : in     vl_logic;
        j_enable_x_qual : in     vl_logic;
        busy_seldr      : in     vl_logic;
        j_com_word4_dat : in     vl_logic_vector(127 downto 0);
        jinstr_cap      : in     vl_logic_vector(7 downto 0);
        jconfig_cap     : in     vl_logic_vector(7 downto 0);
        dsr_out         : in     vl_logic;
        sram_asr_out    : in     vl_logic;
        p8_in           : in     vl_logic_vector(7 downto 0);
        bscan_out       : in     vl_logic;
        isptracy_er1_out: in     vl_logic;
        isptracy_er2_out: in     vl_logic;
        iscan_out       : in     vl_logic_vector(7 downto 0);
        extspi_out      : in     vl_logic
    );
end jtag_register;
