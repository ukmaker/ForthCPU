library verilog;
use verilog.vl_types.all;
entity ser_top is
    port(
        bs4pad_0        : out    vl_logic;
        bs4pad_1        : out    vl_logic;
        bs4refck        : out    vl_logic;
        ck3g4txn2nd     : out    vl_logic;
        ck3g4txp2nd     : out    vl_logic;
        hdoutn0         : out    vl_logic;
        hdoutn1         : out    vl_logic;
        hdoutp0         : out    vl_logic;
        hdoutp1         : out    vl_logic;
        ldr_rx2core     : out    vl_logic_vector(1 downto 0);
        pci_connect0    : out    vl_logic;
        pci_connect1    : out    vl_logic;
        pci_det_done0   : out    vl_logic;
        pci_det_done1   : out    vl_logic;
        plol            : out    vl_logic;
        rck0            : out    vl_logic;
        rck1            : out    vl_logic;
        rd0             : out    vl_logic_vector(9 downto 0);
        rd1             : out    vl_logic_vector(9 downto 0);
        refc2core       : out    vl_logic;
        refck2ndp       : out    vl_logic;
        refck2ndn       : out    vl_logic;
        reg2fpga_out    : out    vl_logic;
        rlol            : out    vl_logic_vector(1 downto 0);
        rx_los          : out    vl_logic_vector(1 downto 0);
        ser_sts_ch0_1   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch0_2   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch0_3   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch1_1   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch1_2   : out    vl_logic_vector(7 downto 0);
        ser_sts_ch1_3   : out    vl_logic_vector(7 downto 0);
        ser_sts_dl_1    : out    vl_logic_vector(7 downto 0);
        sync2ndp        : out    vl_logic;
        sync2ndn        : out    vl_logic;
        tck0            : out    vl_logic;
        tck1            : out    vl_logic;
        tck_aux_full    : out    vl_logic;
        atstn           : inout  vl_logic;
        atstp           : inout  vl_logic;
        vcc             : inout  vl_logic;
        vcca            : inout  vl_logic;
        vcca25          : inout  vl_logic;
        vccarx0         : inout  vl_logic;
        vccarx1         : inout  vl_logic;
        vccatx0         : inout  vl_logic;
        vccatx1         : inout  vl_logic;
        vcchrx0         : inout  vl_logic;
        vcchrx1         : inout  vl_logic;
        vcchtx0         : inout  vl_logic;
        vcchtx1         : inout  vl_logic;
        vss             : inout  vl_logic;
        vssa            : inout  vl_logic;
        vssach0         : inout  vl_logic;
        vssach1         : inout  vl_logic;
        bs2pad_0        : in     vl_logic;
        bs2pad_1        : in     vl_logic;
        cdr_en_bitslip0 : in     vl_logic;
        cdr_en_bitslip1 : in     vl_logic;
        ck3g4txn_nd     : in     vl_logic;
        ck3g4txp_nd     : in     vl_logic;
        ck_core_rx      : in     vl_logic_vector(1 downto 0);
        ck_core_tx      : in     vl_logic;
        hdinn0          : in     vl_logic;
        hdinn1          : in     vl_logic;
        hdinp0          : in     vl_logic;
        hdinp1          : in     vl_logic;
        ib_pwdnb        : in     vl_logic;
        iref_50uconst   : in     vl_logic_vector(1 downto 0);
        iref_50urpoly   : in     vl_logic_vector(1 downto 0);
        ldr_core2tx     : in     vl_logic_vector(1 downto 0);
        macropdb        : in     vl_logic;
        macrorst        : in     vl_logic;
        pci_det_ct0     : in     vl_logic;
        pci_det_ct1     : in     vl_logic;
        pci_det_en0     : in     vl_logic;
        pci_det_en1     : in     vl_logic;
        pci_ei_en0      : in     vl_logic;
        pci_ei_en1      : in     vl_logic;
        pcie_mode       : in     vl_logic_vector(1 downto 0);
        pll_pwdnb       : in     vl_logic;
        pwr_on_rst      : in     vl_logic;
        refck_from_ndp  : in     vl_logic;
        refck_from_ndn  : in     vl_logic;
        refck_pwdnb     : in     vl_logic;
        refclkn         : in     vl_logic;
        refclkp         : in     vl_logic;
        rrst            : in     vl_logic_vector(1 downto 0);
        rx_bs_mode      : in     vl_logic;
        ser_ctl_ch0_1   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_2   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_3   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_4   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_5   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_6   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_7   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_8   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_9   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_10  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_11  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_12  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_13  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch0_14  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_1   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_2   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_3   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_4   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_5   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_6   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_7   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_8   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_9   : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_10  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_11  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_12  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_13  : in     vl_logic_vector(7 downto 0);
        ser_ctl_ch1_14  : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_1    : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_2    : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_3    : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_4    : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_5    : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_6    : in     vl_logic_vector(7 downto 0);
        ser_ctl_dl_7    : in     vl_logic_vector(7 downto 0);
        ser_mem_ch0     : in     vl_logic_vector(87 downto 0);
        ser_mem_ch1     : in     vl_logic_vector(87 downto 0);
        ser_mem_dl      : in     vl_logic_vector(71 downto 0);
        sync_ndp        : in     vl_logic;
        sync_ndn        : in     vl_logic;
        sync_pulse      : in     vl_logic;
        td0             : in     vl_logic_vector(9 downto 0);
        td1             : in     vl_logic_vector(9 downto 0);
        trst            : in     vl_logic;
        tx_bs_mode      : in     vl_logic
    );
end ser_top;
