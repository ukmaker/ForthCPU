library verilog;
use verilog.vl_types.all;
entity pcs_dual_logic is
    port(
        bist_rpt_ch_sel : out    vl_logic;
        bist_rx_clk     : in     vl_logic;
        bist_tx_clk     : in     vl_logic;
        bist_wrst       : in     vl_logic;
        bist_rrst       : in     vl_logic;
        cyawstn         : in     vl_logic;
        ffc_macropdb    : in     vl_logic;
        ffc_sync_toggle : in     vl_logic;
        rstb_txp_1      : in     vl_logic;
        ffs_ls_sync_status: in     vl_logic_vector(1 downto 0);
        mc1_dif_ctl     : in     vl_logic_vector(159 downto 0);
        mc1_ser_ctl_dl  : in     vl_logic_vector(71 downto 0);
        rx_ch           : in     vl_logic_vector(1 downto 0);
        rxr_clk         : in     vl_logic_vector(1 downto 0);
        sciint_10       : in     vl_logic_vector(1 downto 0);
        scirdata_01     : in     vl_logic_vector(7 downto 0);
        sciaddr         : in     vl_logic_vector(5 downto 0);
        scienaux        : in     vl_logic;
        scird           : in     vl_logic;
        sciselaux       : in     vl_logic;
        sciwdata        : in     vl_logic_vector(7 downto 0);
        ser_sts_1_dl_25 : in     vl_logic_vector(7 downto 0);
        tobist_data     : in     vl_logic_vector(9 downto 0);
        reg_load        : in     vl_logic;
        goe_r2          : in     vl_logic;
        goe_load        : in     vl_logic;
        txp_clk1        : in     vl_logic;
        bist_rx_data_sel: out    vl_logic;
        bist_en         : out    vl_logic;
        char_mode       : out    vl_logic;
        fmbist_data     : out    vl_logic_vector(9 downto 0);
        force_int       : out    vl_logic;
        macropdb        : out    vl_logic;
        pcs_ctl_3_dl_02 : out    vl_logic_vector(7 downto 0);
        pcs_ctl_4_dl_03 : out    vl_logic_vector(7 downto 0);
        rst_ctl_1_dl_10 : out    vl_logic_vector(7 downto 0);
        sciint          : out    vl_logic;
        scirdata        : out    vl_logic_vector(7 downto 0);
        ser_ctl_1_dl_0a : out    vl_logic_vector(7 downto 0);
        ser_ctl_2_dl_0b : out    vl_logic_vector(7 downto 0);
        ser_ctl_3_dl_0c : out    vl_logic_vector(7 downto 0);
        ser_ctl_4_dl_0d : out    vl_logic_vector(7 downto 0);
        ser_ctl_5_dl_0e : out    vl_logic_vector(7 downto 0);
        ser_ctl_6_dl_12 : out    vl_logic_vector(7 downto 0);
        ser_ctl_7_dl_13 : out    vl_logic_vector(7 downto 0);
        sync_pulse      : out    vl_logic;
        xge_mode        : out    vl_logic;
        ser_mem_dl      : out    vl_logic_vector(71 downto 0)
    );
end pcs_dual_logic;
