library verilog;
use verilog.vl_types.all;
entity EFB is
    generic(
        EFB_I2C1        : string  := "DISABLED";
        EFB_I2C2        : string  := "DISABLED";
        EFB_SPI         : string  := "DISABLED";
        EFB_TC          : string  := "DISABLED";
        EFB_TC_PORTMODE : string  := "NO_WB";
        EFB_UFM         : string  := "DISABLED";
        EFB_WB_CLK_FREQ : string  := "50.0";
        DEV_DENSITY     : string  := "1200L";
        UFM_INIT_PAGES  : integer := 0;
        UFM_INIT_START_PAGE: integer := 0;
        UFM_INIT_ALL_ZEROS: string  := "ENABLED";
        UFM_INIT_FILE_NAME: string  := "NONE";
        UFM_INIT_FILE_FORMAT: string  := "HEX";
        I2C1_ADDRESSING : string  := "7BIT";
        I2C2_ADDRESSING : string  := "7BIT";
        I2C1_SLAVE_ADDR : string  := "0b1000001";
        I2C2_SLAVE_ADDR : string  := "0b1000010";
        I2C1_BUS_PERF   : string  := "100kHz";
        I2C2_BUS_PERF   : string  := "100kHz";
        I2C1_CLK_DIVIDER: integer := 1;
        I2C2_CLK_DIVIDER: integer := 1;
        I2C1_GEN_CALL   : string  := "DISABLED";
        I2C2_GEN_CALL   : string  := "DISABLED";
        I2C1_WAKEUP     : string  := "DISABLED";
        I2C2_WAKEUP     : string  := "DISABLED";
        SPI_MODE        : string  := "SLAVE";
        SPI_CLK_DIVIDER : integer := 1;
        SPI_LSB_FIRST   : string  := "DISABLED";
        SPI_CLK_INV     : string  := "DISABLED";
        SPI_PHASE_ADJ   : string  := "DISABLED";
        SPI_SLAVE_HANDSHAKE: string  := "DISABLED";
        SPI_INTR_TXRDY  : string  := "DISABLED";
        SPI_INTR_RXRDY  : string  := "DISABLED";
        SPI_INTR_TXOVR  : string  := "DISABLED";
        SPI_INTR_RXOVR  : string  := "DISABLED";
        SPI_WAKEUP      : string  := "DISABLED";
        TC_MODE         : string  := "CTCM";
        TC_SCLK_SEL     : string  := "PCLOCK";
        TC_CCLK_SEL     : integer := 1;
        GSR             : string  := "ENABLED";
        TC_TOP_SET      : integer := 65535;
        TC_OCR_SET      : integer := 32767;
        TC_OC_MODE      : string  := "TOGGLE";
        TC_RESETN       : string  := "ENABLED";
        TC_TOP_SEL      : string  := "ON";
        TC_OV_INT       : string  := "OFF";
        TC_OCR_INT      : string  := "OFF";
        TC_ICR_INT      : string  := "OFF";
        TC_OVERFLOW     : string  := "ENABLED";
        TC_ICAPTURE     : string  := "DISABLED"
    );
    port(
        WBCLKI          : in     vl_logic;
        WBRSTI          : in     vl_logic;
        WBCYCI          : in     vl_logic;
        WBSTBI          : in     vl_logic;
        WBWEI           : in     vl_logic;
        WBADRI7         : in     vl_logic;
        WBADRI6         : in     vl_logic;
        WBADRI5         : in     vl_logic;
        WBADRI4         : in     vl_logic;
        WBADRI3         : in     vl_logic;
        WBADRI2         : in     vl_logic;
        WBADRI1         : in     vl_logic;
        WBADRI0         : in     vl_logic;
        WBDATI7         : in     vl_logic;
        WBDATI6         : in     vl_logic;
        WBDATI5         : in     vl_logic;
        WBDATI4         : in     vl_logic;
        WBDATI3         : in     vl_logic;
        WBDATI2         : in     vl_logic;
        WBDATI1         : in     vl_logic;
        WBDATI0         : in     vl_logic;
        PLL0DATI7       : in     vl_logic;
        PLL0DATI6       : in     vl_logic;
        PLL0DATI5       : in     vl_logic;
        PLL0DATI4       : in     vl_logic;
        PLL0DATI3       : in     vl_logic;
        PLL0DATI2       : in     vl_logic;
        PLL0DATI1       : in     vl_logic;
        PLL0DATI0       : in     vl_logic;
        PLL0ACKI        : in     vl_logic;
        PLL1DATI7       : in     vl_logic;
        PLL1DATI6       : in     vl_logic;
        PLL1DATI5       : in     vl_logic;
        PLL1DATI4       : in     vl_logic;
        PLL1DATI3       : in     vl_logic;
        PLL1DATI2       : in     vl_logic;
        PLL1DATI1       : in     vl_logic;
        PLL1DATI0       : in     vl_logic;
        PLL1ACKI        : in     vl_logic;
        I2C1SCLI        : in     vl_logic;
        I2C1SDAI        : in     vl_logic;
        I2C2SCLI        : in     vl_logic;
        I2C2SDAI        : in     vl_logic;
        SPISCKI         : in     vl_logic;
        SPIMISOI        : in     vl_logic;
        SPIMOSII        : in     vl_logic;
        SPISCSN         : in     vl_logic;
        TCCLKI          : in     vl_logic;
        TCRSTN          : in     vl_logic;
        TCIC            : in     vl_logic;
        UFMSN           : in     vl_logic;
        WBDATO7         : out    vl_logic;
        WBDATO6         : out    vl_logic;
        WBDATO5         : out    vl_logic;
        WBDATO4         : out    vl_logic;
        WBDATO3         : out    vl_logic;
        WBDATO2         : out    vl_logic;
        WBDATO1         : out    vl_logic;
        WBDATO0         : out    vl_logic;
        WBACKO          : out    vl_logic;
        PLLCLKO         : out    vl_logic;
        PLLRSTO         : out    vl_logic;
        PLL0STBO        : out    vl_logic;
        PLL1STBO        : out    vl_logic;
        PLLWEO          : out    vl_logic;
        PLLADRO4        : out    vl_logic;
        PLLADRO3        : out    vl_logic;
        PLLADRO2        : out    vl_logic;
        PLLADRO1        : out    vl_logic;
        PLLADRO0        : out    vl_logic;
        PLLDATO7        : out    vl_logic;
        PLLDATO6        : out    vl_logic;
        PLLDATO5        : out    vl_logic;
        PLLDATO4        : out    vl_logic;
        PLLDATO3        : out    vl_logic;
        PLLDATO2        : out    vl_logic;
        PLLDATO1        : out    vl_logic;
        PLLDATO0        : out    vl_logic;
        WBCUFMIRQ       : out    vl_logic;
        I2C1SCLO        : out    vl_logic;
        I2C1SCLOEN      : out    vl_logic;
        I2C1SDAO        : out    vl_logic;
        I2C1SDAOEN      : out    vl_logic;
        I2C2SCLO        : out    vl_logic;
        I2C2SCLOEN      : out    vl_logic;
        I2C2SDAO        : out    vl_logic;
        I2C2SDAOEN      : out    vl_logic;
        I2C1IRQO        : out    vl_logic;
        I2C2IRQO        : out    vl_logic;
        SPISCKO         : out    vl_logic;
        SPISCKEN        : out    vl_logic;
        SPIMISOO        : out    vl_logic;
        SPIMISOEN       : out    vl_logic;
        SPIMOSIO        : out    vl_logic;
        SPIMOSIEN       : out    vl_logic;
        SPIMCSN0        : out    vl_logic;
        SPIMCSN1        : out    vl_logic;
        SPIMCSN2        : out    vl_logic;
        SPIMCSN3        : out    vl_logic;
        SPIMCSN4        : out    vl_logic;
        SPIMCSN5        : out    vl_logic;
        SPIMCSN6        : out    vl_logic;
        SPIMCSN7        : out    vl_logic;
        SPICSNEN        : out    vl_logic;
        SPIIRQO         : out    vl_logic;
        TCINT           : out    vl_logic;
        TCOC            : out    vl_logic;
        CFGWAKE         : out    vl_logic;
        CFGSTDBY        : out    vl_logic
    );
end EFB;
