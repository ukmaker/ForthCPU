library verilog;
use verilog.vl_types.all;
entity delc1x2v1s is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end delc1x2v1s;
