library verilog;
use verilog.vl_types.all;
entity spare_gate_efb_1 is
    port(
        signal_in       : in     vl_logic
    );
end spare_gate_efb_1;
