library verilog;
use verilog.vl_types.all;
entity BUFX4 is
    port(
        z               : out    vl_logic;
        a               : in     vl_logic
    );
end BUFX4;
