library verilog;
use verilog.vl_types.all;
entity njtag_register is
    port(
        njcommand       : out    vl_logic_vector(7 downto 0);
        njconfig_dat    : out    vl_logic_vector(3 downto 0);
        njsector_dat    : out    vl_logic_vector(7 downto 0);
        njbuf128_dat    : out    vl_logic_vector(127 downto 0);
        njcom_out       : out    vl_logic_vector(7 downto 0);
        nj_load_op2     : out    vl_logic;
        nj_load_op3     : out    vl_logic;
        nj_operand1     : out    vl_logic_vector(7 downto 0);
        nj_operand2     : out    vl_logic_vector(7 downto 0);
        nj_operand3     : out    vl_logic_vector(7 downto 0);
        cmd_noop        : out    vl_logic;
        nj_check_crc_en : out    vl_logic;
        nj_rcv_rd_cmd   : out    vl_logic;
        nj_dsr_data     : out    vl_logic_vector(7 downto 0);
        nj_jump_param   : out    vl_logic_vector(31 downto 0);
        nj_csel_param   : out    vl_logic_vector(7 downto 0);
        njpspi_ctrl     : out    vl_logic_vector(15 downto 0);
        njpcs_addr_dat  : out    vl_logic_vector(14 downto 0);
        por             : in     vl_logic;
        smclk           : in     vl_logic;
        ref_launch      : in     vl_logic;
        nj_rst_sync     : in     vl_logic;
        njcmd_dec       : in     vl_logic;
        njcmd_inf1      : in     vl_logic;
        njcmd_inf2      : in     vl_logic;
        njcmd_inf3      : in     vl_logic;
        nj_exec_a       : in     vl_logic;
        nj_exec_b       : in     vl_logic;
        nj_exec_f       : in     vl_logic;
        njtag_din       : in     vl_logic_vector(7 downto 0);
        njtag_run       : in     vl_logic;
        com_shift_en    : in     vl_logic;
        ctrl_wkup_tran  : in     vl_logic;
        njsel_cfg       : in     vl_logic;
        njsel_sec       : in     vl_logic;
        njsel_com       : in     vl_logic;
        njsel_extspi    : in     vl_logic;
        njcap_com_word4_norm: in     vl_logic;
        njcap_com_word4_slow: in     vl_logic;
        njshf_com_byte1 : in     vl_logic;
        njshf_com_byte2 : in     vl_logic;
        njshf_com_byte4 : in     vl_logic;
        njshf_com_byte8 : in     vl_logic;
        njshf_com_byte9 : in     vl_logic;
        njshf_com_word4 : in     vl_logic;
        nj_enable_qual  : in     vl_logic;
        nj_enable_x_qual: in     vl_logic;
        lsc_pcs_rw_c    : in     vl_logic;
        nj_cmd_prog_dsr : in     vl_logic;
        nj_cmd_read_dat : in     vl_logic;
        nj_cmd_read     : in     vl_logic;
        nj_com_word4_dat: in     vl_logic_vector(127 downto 0);
        njtag_slow_response: in     vl_logic
    );
end njtag_register;
