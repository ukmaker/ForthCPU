library verilog;
use verilog.vl_types.all;
entity ser_rx_top is
    port(
        bsout_rx        : out    vl_logic;
        dco_calib_done  : out    vl_logic;
        dco_calib_err   : out    vl_logic;
        dco_facq_done   : out    vl_logic;
        dco_facq_err    : out    vl_logic;
        dco_status      : out    vl_logic_vector(15 downto 0);
        rck             : out    vl_logic;
        rd              : out    vl_logic_vector(9 downto 0);
        rlol            : out    vl_logic;
        rx_hstest1      : out    vl_logic;
        rx_los          : out    vl_logic;
        slb_dn          : out    vl_logic;
        slb_dp          : out    vl_logic;
        slb_r2t         : out    vl_logic;
        slb_r2tb        : out    vl_logic;
        i50u4dco_const  : inout  vl_logic_vector(1 downto 0);
        i50u4leq_const  : inout  vl_logic_vector(1 downto 0);
        i50u4leq_poly   : inout  vl_logic_vector(1 downto 0);
        i50u4pd_poly    : inout  vl_logic_vector(1 downto 0);
        i50u4rxbs_poly  : inout  vl_logic;
        vcc             : inout  vl_logic;
        vcca25          : inout  vl_logic;
        vccarx          : inout  vl_logic;
        vcchrx          : inout  vl_logic;
        vss             : inout  vl_logic;
        vssarx          : inout  vl_logic;
        vssarxs         : inout  vl_logic;
        atsten          : in     vl_logic;
        auto_calib_en   : in     vl_logic;
        auto_facq_en    : in     vl_logic;
        band_calib_mode : in     vl_logic;
        band_threshold  : in     vl_logic_vector(5 downto 0);
        bs_mode         : in     vl_logic;
        bus8bit_sel     : in     vl_logic;
        calib_ck_mode   : in     vl_logic;
        calib_time_sel  : in     vl_logic_vector(1 downto 0);
        cdr_dlock       : in     vl_logic;
        cdr_en_bitslip  : in     vl_logic;
        cdr_lol_set     : in     vl_logic_vector(1 downto 0);
        ck_core_rx      : in     vl_logic;
        dac_bdavoid_enb : in     vl_logic;
        dco_calib_rst   : in     vl_logic;
        dco_facq_rst    : in     vl_logic;
        div11en_rx      : in     vl_logic;
        dnlb            : in     vl_logic;
        dplb            : in     vl_logic;
        en_recalib      : in     vl_logic;
        fc2dco_dloop    : in     vl_logic;
        fc2dco_floop    : in     vl_logic;
        hdinn           : in     vl_logic;
        hdinp           : in     vl_logic;
        lb_ctl          : in     vl_logic_vector(3 downto 0);
        leq_offset_sel  : in     vl_logic;
        leq_offset_trim : in     vl_logic_vector(2 downto 0);
        pd_iset         : in     vl_logic_vector(1 downto 0);
        pden_sel        : in     vl_logic;
        rate_mode_rx    : in     vl_logic;
        rate_sel        : in     vl_logic_vector(3 downto 0);
        rcv_dcc_en      : in     vl_logic;
        refck25x        : in     vl_logic;
        refck_mode      : in     vl_logic_vector(1 downto 0);
        refck_modeo     : in     vl_logic_vector(1 downto 0);
        reg_band_offset : in     vl_logic_vector(3 downto 0);
        reg_band_sel    : in     vl_logic_vector(5 downto 0);
        reg_idac_en     : in     vl_logic;
        reg_idac_sel    : in     vl_logic_vector(9 downto 0);
        req_en          : in     vl_logic;
        req_iset        : in     vl_logic_vector(2 downto 0);
        req_lvl_set     : in     vl_logic_vector(1 downto 0);
        reset_vcc       : in     vl_logic;
        resetb          : in     vl_logic;
        rlos_sel        : in     vl_logic;
        rlos_vcc        : in     vl_logic;
        rpwdnb          : in     vl_logic;
        rrst            : in     vl_logic;
        rterm_rx        : in     vl_logic_vector(3 downto 0);
        rx_dco_ck_div   : in     vl_logic_vector(2 downto 0);
        rx_ldr_sel      : in     vl_logic;
        rx_los_ceq      : in     vl_logic_vector(1 downto 0);
        rx_los_en       : in     vl_logic;
        rx_los_hyst_en  : in     vl_logic;
        rx_los_lvl      : in     vl_logic_vector(2 downto 0);
        rx_refck_local  : in     vl_logic;
        rx_refck_sel    : in     vl_logic;
        rx_spare_inb    : in     vl_logic_vector(7 downto 0);
        rx_spare_inc    : in     vl_logic_vector(7 downto 0);
        rxin_cm         : in     vl_logic_vector(1 downto 0);
        rxterm_cm       : in     vl_logic_vector(1 downto 0);
        ser_mem         : in     vl_logic_vector(43 downto 0)
    );
end ser_rx_top;
