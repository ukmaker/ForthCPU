library verilog;
use verilog.vl_types.all;
entity model_top_reno is
    port(
        ana_rst_b       : out    vl_logic;
        ascclk_oeb      : out    vl_logic;
        ascclk_out      : out    vl_logic;
        bpz             : out    vl_logic_vector(1 downto 0);
        cfg_hvout       : out    vl_logic_vector(31 downto 0);
        cfg_im          : out    vl_logic_vector(30 downto 0);
        clk_loss_off    : out    vl_logic;
        dac_resetb      : out    vl_logic;
        dacin           : out    vl_logic_vector(7 downto 0);
        dtpi_en         : out    vl_logic;
        dtpo            : out    vl_logic;
        dtpo_en         : out    vl_logic;
        gpio_oeb        : out    vl_logic_vector(10 downto 1);
        gpio_out        : out    vl_logic_vector(10 downto 1);
        gpio_pldn_en    : out    vl_logic_vector(10 downto 1);
        hvout_data      : out    vl_logic_vector(4 downto 1);
        i2cdet_clk      : out    vl_logic;
        i2cdet_resetb   : out    vl_logic;
        i2cdet_tapsel   : out    vl_logic_vector(2 downto 0);
        im_hc_en        : out    vl_logic_vector(1 downto 0);
        ldmshdw         : out    vl_logic;
        ldshdwreg       : out    vl_logic;
        ldsshdw         : out    vl_logic;
        mclk            : out    vl_logic;
        mfg_abg         : out    vl_logic_vector(12 downto 0);
        mfg_abg_enb     : out    vl_logic;
        mfg_adc_enb     : out    vl_logic;
        mfg_dac         : out    vl_logic_vector(4 downto 0);
        mfg_dac_enb     : out    vl_logic;
        mfg_en_atp1     : out    vl_logic;
        mfg_en_atp2     : out    vl_logic;
        mfg_en_dtpi     : out    vl_logic;
        mfg_en_dtpo     : out    vl_logic;
        mfg_en_matp1    : out    vl_logic;
        mfg_en_matp2    : out    vl_logic;
        mfg_hvblk_dis   : out    vl_logic;
        mfg_i2cdet      : out    vl_logic;
        mfg_im          : out    vl_logic_vector(6 downto 0);
        mfg_osc_vref    : out    vl_logic;
        mfg_sar_m_en    : out    vl_logic;
        mfg_sar_p_en    : out    vl_logic;
        mfg_sp          : out    vl_logic_vector(3 downto 0);
        mfg_tm          : out    vl_logic_vector(7 downto 0);
        mfg_vm          : out    vl_logic;
        mfg_vmon_bypass : out    vl_logic;
        mfg_vmon_enb    : out    vl_logic;
        por_off         : out    vl_logic;
        rdat            : out    vl_logic;
        rdat_oeb        : out    vl_logic;
        rdshdw          : out    vl_logic;
        reset_in_b      : out    vl_logic;
        resetb_out_pin  : out    vl_logic;
        rst_abg_b       : out    vl_logic;
        rst_clk_gen_b   : out    vl_logic;
        rst_osc_b       : out    vl_logic;
        rst_osc_tmr_b   : out    vl_logic;
        safestate       : out    vl_logic;
        sar_atten       : out    vl_logic;
        sar_muxsel      : out    vl_logic_vector(3 downto 0);
        sar_socb        : out    vl_logic;
        sda_out         : out    vl_logic;
        tm_adc_clk      : out    vl_logic;
        tm_adc_resetb   : out    vl_logic;
        tm_beta_done    : out    vl_logic;
        tm_beta_en      : out    vl_logic;
        tm_betabits     : out    vl_logic_vector(5 downto 0);
        tm_chansel      : out    vl_logic_vector(2 downto 0);
        tm_demout       : out    vl_logic;
        tm_demratio     : out    vl_logic_vector(15 downto 0);
        tm_porkchop     : out    vl_logic;
        tm_single_e     : out    vl_logic;
        trim_bg_buff    : out    vl_logic_vector(27 downto 0);
        trim_dac        : out    vl_logic_vector(3 downto 0);
        trim_osc        : out    vl_logic_vector(3 downto 0);
        trim_osc_vref   : out    vl_logic_vector(2 downto 0);
        trim_se_deriv   : out    vl_logic;
        trim_sp_bg      : out    vl_logic_vector(4 downto 0);
        trim_tm         : out    vl_logic;
        trimoutenable   : out    vl_logic_vector(3 downto 0);
        vdbg            : out    vl_logic;
        vhi             : out    vl_logic;
        vmon_hc_en      : out    vl_logic_vector(1 downto 0);
        cfg_vm          : inout  vl_logic_vector(7 downto 0);
        iabias_25u      : inout  vl_logic;
        ihvout0_n5u     : inout  vl_logic;
        ihvout1_n5u     : inout  vl_logic;
        ihvout2_n5u     : inout  vl_logic;
        ihvout3_n5u     : inout  vl_logic;
        ii2c_25u        : inout  vl_logic;
        ioa_25u         : inout  vl_logic;
        iosc_25u        : inout  vl_logic;
        irefpad_bot10u  : inout  vl_logic;
        irefpad_top10u  : inout  vl_logic;
        matp1           : inout  vl_logic;
        matp2           : inout  vl_logic;
        vddd            : inout  vl_logic;
        vpp             : inout  vl_logic;
        vssd            : inout  vl_logic;
        bg_caldone      : in     vl_logic;
        dac_chan        : in     vl_logic_vector(2 downto 0);
        dac_init        : in     vl_logic;
        dac_ready       : in     vl_logic;
        dtpi            : in     vl_logic;
        fsafeb          : in     vl_logic;
        gpio_in         : in     vl_logic_vector(10 downto 1);
        hvblock         : in     vl_logic;
        i2cdet_compout  : in     vl_logic;
        im_fcout        : in     vl_logic;
        im_gf_a         : in     vl_logic;
        im_gf_b         : in     vl_logic;
        imhv_fcout      : in     vl_logic;
        imhv_gf_a       : in     vl_logic;
        imhv_gf_b       : in     vl_logic;
        mclkout         : in     vl_logic;
        por_n           : in     vl_logic;
        resetb_in_pin   : in     vl_logic;
        sar_data        : in     vl_logic_vector(9 downto 0);
        sar_done        : in     vl_logic;
        scl_in          : in     vl_logic;
        sda_in          : in     vl_logic;
        sync_hvblk      : in     vl_logic;
        tm_betacomp     : in     vl_logic;
        tm_modout       : in     vl_logic;
        v2p1            : in     vl_logic;
        vmon_odd        : in     vl_logic;
        vmona           : in     vl_logic_vector(10 downto 1);
        vmonb           : in     vl_logic_vector(10 downto 1);
        wdat            : in     vl_logic;
        tmon_1a         : in     vl_logic;
        tmon_1b         : in     vl_logic;
        tmon_2a         : in     vl_logic;
        tmon_2b         : in     vl_logic;
        tmonint_1a      : in     vl_logic;
        tmonint_1b      : in     vl_logic;
        wrclk_in        : in     vl_logic;
        wrclk_lost      : in     vl_logic
    );
end model_top_reno;
