library verilog;
use verilog.vl_types.all;
entity DCUA is
    generic(
        D_MACROPDB      : string  := "DONTCARE";
        D_IB_PWDNB      : string  := "DONTCARE";
        D_XGE_MODE      : string  := "DONTCARE";
        D_LOW_MARK      : string  := "DONTCARE";
        D_HIGH_MARK     : string  := "DONTCARE";
        D_BUS8BIT_SEL   : string  := "DONTCARE";
        D_CDR_LOL_SET   : string  := "DONTCARE";
        D_BITCLK_LOCAL_EN: string  := "DONTCARE";
        D_BITCLK_ND_EN  : string  := "DONTCARE";
        D_BITCLK_FROM_ND_EN: string  := "DONTCARE";
        D_SYNC_LOCAL_EN : string  := "DONTCARE";
        D_SYNC_ND_EN    : string  := "DONTCARE";
        CH0_UC_MODE     : string  := "DONTCARE";
        CH1_UC_MODE     : string  := "DONTCARE";
        CH0_PCIE_MODE   : string  := "DONTCARE";
        CH1_PCIE_MODE   : string  := "DONTCARE";
        CH0_RIO_MODE    : string  := "DONTCARE";
        CH1_RIO_MODE    : string  := "DONTCARE";
        CH0_WA_MODE     : string  := "DONTCARE";
        CH1_WA_MODE     : string  := "DONTCARE";
        CH0_INVERT_RX   : string  := "DONTCARE";
        CH1_INVERT_RX   : string  := "DONTCARE";
        CH0_INVERT_TX   : string  := "DONTCARE";
        CH1_INVERT_TX   : string  := "DONTCARE";
        CH0_PRBS_SELECTION: string  := "DONTCARE";
        CH1_PRBS_SELECTION: string  := "DONTCARE";
        CH0_GE_AN_ENABLE: string  := "DONTCARE";
        CH1_GE_AN_ENABLE: string  := "DONTCARE";
        CH0_PRBS_LOCK   : string  := "DONTCARE";
        CH1_PRBS_LOCK   : string  := "DONTCARE";
        CH0_PRBS_ENABLE : string  := "DONTCARE";
        CH1_PRBS_ENABLE : string  := "DONTCARE";
        CH0_ENABLE_CG_ALIGN: string  := "DONTCARE";
        CH1_ENABLE_CG_ALIGN: string  := "DONTCARE";
        CH0_TX_GEAR_MODE: string  := "DONTCARE";
        CH1_TX_GEAR_MODE: string  := "DONTCARE";
        CH0_RX_GEAR_MODE: string  := "DONTCARE";
        CH1_RX_GEAR_MODE: string  := "DONTCARE";
        CH0_PCS_DET_TIME_SEL: string  := "DONTCARE";
        CH1_PCS_DET_TIME_SEL: string  := "DONTCARE";
        CH0_PCIE_EI_EN  : string  := "DONTCARE";
        CH1_PCIE_EI_EN  : string  := "DONTCARE";
        CH0_TX_GEAR_BYPASS: string  := "DONTCARE";
        CH1_TX_GEAR_BYPASS: string  := "DONTCARE";
        CH0_ENC_BYPASS  : string  := "DONTCARE";
        CH1_ENC_BYPASS  : string  := "DONTCARE";
        CH0_SB_BYPASS   : string  := "DONTCARE";
        CH1_SB_BYPASS   : string  := "DONTCARE";
        CH0_RX_SB_BYPASS: string  := "DONTCARE";
        CH1_RX_SB_BYPASS: string  := "DONTCARE";
        CH0_WA_BYPASS   : string  := "DONTCARE";
        CH1_WA_BYPASS   : string  := "DONTCARE";
        CH0_DEC_BYPASS  : string  := "DONTCARE";
        CH1_DEC_BYPASS  : string  := "DONTCARE";
        CH0_CTC_BYPASS  : string  := "DONTCARE";
        CH1_CTC_BYPASS  : string  := "DONTCARE";
        CH0_RX_GEAR_BYPASS: string  := "DONTCARE";
        CH1_RX_GEAR_BYPASS: string  := "DONTCARE";
        CH0_LSM_DISABLE : string  := "DONTCARE";
        CH1_LSM_DISABLE : string  := "DONTCARE";
        CH0_MATCH_2_ENABLE: string  := "DONTCARE";
        CH1_MATCH_2_ENABLE: string  := "DONTCARE";
        CH0_MATCH_4_ENABLE: string  := "DONTCARE";
        CH1_MATCH_4_ENABLE: string  := "DONTCARE";
        CH0_MIN_IPG_CNT : string  := "DONTCARE";
        CH1_MIN_IPG_CNT : string  := "DONTCARE";
        CH0_CC_MATCH_1  : string  := "DONTCARE";
        CH1_CC_MATCH_1  : string  := "DONTCARE";
        CH0_CC_MATCH_2  : string  := "DONTCARE";
        CH1_CC_MATCH_2  : string  := "DONTCARE";
        CH0_CC_MATCH_3  : string  := "DONTCARE";
        CH1_CC_MATCH_3  : string  := "DONTCARE";
        CH0_CC_MATCH_4  : string  := "DONTCARE";
        CH1_CC_MATCH_4  : string  := "DONTCARE";
        CH0_UDF_COMMA_MASK: string  := "DONTCARE";
        CH1_UDF_COMMA_MASK: string  := "DONTCARE";
        CH0_UDF_COMMA_A : string  := "DONTCARE";
        CH1_UDF_COMMA_A : string  := "DONTCARE";
        CH0_UDF_COMMA_B : string  := "DONTCARE";
        CH1_UDF_COMMA_B : string  := "DONTCARE";
        CH0_RX_DCO_CK_DIV: string  := "DONTCARE";
        CH1_RX_DCO_CK_DIV: string  := "DONTCARE";
        CH0_RCV_DCC_EN  : string  := "DONTCARE";
        CH1_RCV_DCC_EN  : string  := "DONTCARE";
        CH0_REQ_LVL_SET : string  := "DONTCARE";
        CH1_REQ_LVL_SET : string  := "DONTCARE";
        CH0_REQ_EN      : string  := "DONTCARE";
        CH1_REQ_EN      : string  := "DONTCARE";
        CH0_RTERM_RX    : string  := "DONTCARE";
        CH1_RTERM_RX    : string  := "DONTCARE";
        CH0_PDEN_SEL    : string  := "DONTCARE";
        CH1_PDEN_SEL    : string  := "DONTCARE";
        CH0_TPWDNB      : string  := "DONTCARE";
        CH1_TPWDNB      : string  := "DONTCARE";
        CH0_RATE_MODE_TX: string  := "DONTCARE";
        CH1_RATE_MODE_TX: string  := "DONTCARE";
        CH0_RTERM_TX    : string  := "DONTCARE";
        CH1_RTERM_TX    : string  := "DONTCARE";
        CH0_TX_CM_SEL   : string  := "DONTCARE";
        CH1_TX_CM_SEL   : string  := "DONTCARE";
        CH0_TDRV_PRE_EN : string  := "DONTCARE";
        CH1_TDRV_PRE_EN : string  := "DONTCARE";
        CH0_TDRV_SLICE0_SEL: string  := "DONTCARE";
        CH1_TDRV_SLICE0_SEL: string  := "DONTCARE";
        CH0_TDRV_SLICE1_SEL: string  := "DONTCARE";
        CH1_TDRV_SLICE1_SEL: string  := "DONTCARE";
        CH0_TDRV_SLICE2_SEL: string  := "DONTCARE";
        CH1_TDRV_SLICE2_SEL: string  := "DONTCARE";
        CH0_TDRV_SLICE3_SEL: string  := "DONTCARE";
        CH1_TDRV_SLICE3_SEL: string  := "DONTCARE";
        CH0_TDRV_SLICE4_SEL: string  := "DONTCARE";
        CH1_TDRV_SLICE4_SEL: string  := "DONTCARE";
        CH0_TDRV_SLICE5_SEL: string  := "DONTCARE";
        CH1_TDRV_SLICE5_SEL: string  := "DONTCARE";
        CH0_TDRV_SLICE0_CUR: string  := "DONTCARE";
        CH1_TDRV_SLICE0_CUR: string  := "DONTCARE";
        CH0_TDRV_SLICE1_CUR: string  := "DONTCARE";
        CH1_TDRV_SLICE1_CUR: string  := "DONTCARE";
        CH0_TDRV_SLICE2_CUR: string  := "DONTCARE";
        CH1_TDRV_SLICE2_CUR: string  := "DONTCARE";
        CH0_TDRV_SLICE3_CUR: string  := "DONTCARE";
        CH1_TDRV_SLICE3_CUR: string  := "DONTCARE";
        CH0_TDRV_SLICE4_CUR: string  := "DONTCARE";
        CH1_TDRV_SLICE4_CUR: string  := "DONTCARE";
        CH0_TDRV_SLICE5_CUR: string  := "DONTCARE";
        CH1_TDRV_SLICE5_CUR: string  := "DONTCARE";
        CH0_TDRV_DAT_SEL: string  := "DONTCARE";
        CH1_TDRV_DAT_SEL: string  := "DONTCARE";
        CH0_TX_DIV11_SEL: string  := "DONTCARE";
        CH1_TX_DIV11_SEL: string  := "DONTCARE";
        CH0_RPWDNB      : string  := "DONTCARE";
        CH1_RPWDNB      : string  := "DONTCARE";
        CH0_RATE_MODE_RX: string  := "DONTCARE";
        CH1_RATE_MODE_RX: string  := "DONTCARE";
        CH0_RLOS_SEL    : string  := "DONTCARE";
        CH1_RLOS_SEL    : string  := "DONTCARE";
        CH0_RX_LOS_LVL  : string  := "DONTCARE";
        CH1_RX_LOS_LVL  : string  := "DONTCARE";
        CH0_RX_LOS_CEQ  : string  := "DONTCARE";
        CH1_RX_LOS_CEQ  : string  := "DONTCARE";
        CH0_RX_LOS_HYST_EN: string  := "DONTCARE";
        CH1_RX_LOS_HYST_EN: string  := "DONTCARE";
        CH0_RX_LOS_EN   : string  := "DONTCARE";
        CH1_RX_LOS_EN   : string  := "DONTCARE";
        CH0_RX_DIV11_SEL: string  := "DONTCARE";
        CH1_RX_DIV11_SEL: string  := "DONTCARE";
        CH0_SEL_SD_RX_CLK: string  := "DONTCARE";
        CH1_SEL_SD_RX_CLK: string  := "DONTCARE";
        CH0_FF_RX_H_CLK_EN: string  := "DONTCARE";
        CH1_FF_RX_H_CLK_EN: string  := "DONTCARE";
        CH0_FF_RX_F_CLK_DIS: string  := "DONTCARE";
        CH1_FF_RX_F_CLK_DIS: string  := "DONTCARE";
        CH0_FF_TX_H_CLK_EN: string  := "DONTCARE";
        CH1_FF_TX_H_CLK_EN: string  := "DONTCARE";
        CH0_FF_TX_F_CLK_DIS: string  := "DONTCARE";
        CH1_FF_TX_F_CLK_DIS: string  := "DONTCARE";
        CH0_RX_RATE_SEL : string  := "DONTCARE";
        CH1_RX_RATE_SEL : string  := "DONTCARE";
        CH0_TDRV_POST_EN: string  := "DONTCARE";
        CH1_TDRV_POST_EN: string  := "DONTCARE";
        CH0_TX_POST_SIGN: string  := "DONTCARE";
        CH1_TX_POST_SIGN: string  := "DONTCARE";
        CH0_TX_PRE_SIGN : string  := "DONTCARE";
        CH1_TX_PRE_SIGN : string  := "DONTCARE";
        CH0_RXTERM_CM   : string  := "DONTCARE";
        CH1_RXTERM_CM   : string  := "DONTCARE";
        CH0_RXIN_CM     : string  := "DONTCARE";
        CH1_RXIN_CM     : string  := "DONTCARE";
        CH0_LEQ_OFFSET_SEL: string  := "DONTCARE";
        CH1_LEQ_OFFSET_SEL: string  := "DONTCARE";
        CH0_LEQ_OFFSET_TRIM: string  := "DONTCARE";
        CH1_LEQ_OFFSET_TRIM: string  := "DONTCARE";
        CH0_LDR_RX2CORE_SEL: string  := "DONTCARE";
        CH1_LDR_RX2CORE_SEL: string  := "DONTCARE";
        CH0_LDR_CORE2TX_SEL: string  := "DONTCARE";
        CH1_LDR_CORE2TX_SEL: string  := "DONTCARE";
        D_TX_MAX_RATE   : string  := "DONTCARE";
        CH0_CDR_MAX_RATE: string  := "DONTCARE";
        CH1_CDR_MAX_RATE: string  := "DONTCARE";
        CH0_TXAMPLITUDE : string  := "DONTCARE";
        CH1_TXAMPLITUDE : string  := "DONTCARE";
        CH0_TXDEPRE     : string  := "DONTCARE";
        CH1_TXDEPRE     : string  := "DONTCARE";
        CH0_TXDEPOST    : string  := "DONTCARE";
        CH1_TXDEPOST    : string  := "DONTCARE";
        CH0_PROTOCOL    : string  := "DONTCARE";
        CH1_PROTOCOL    : string  := "DONTCARE";
        D_ISETLOS       : string  := "DONTCARE";
        D_SETIRPOLY_AUX : string  := "DONTCARE";
        D_SETICONST_AUX : string  := "DONTCARE";
        D_SETIRPOLY_CH  : string  := "DONTCARE";
        D_SETICONST_CH  : string  := "DONTCARE";
        D_REQ_ISET      : string  := "DONTCARE";
        D_PD_ISET       : string  := "DONTCARE";
        D_DCO_CALIB_TIME_SEL: string  := "DONTCARE";
        CH0_DCOCTLGI    : string  := "DONTCARE";
        CH1_DCOCTLGI    : string  := "DONTCARE";
        CH0_DCOATDDLY   : string  := "DONTCARE";
        CH1_DCOATDDLY   : string  := "DONTCARE";
        CH0_DCOATDCFG   : string  := "DONTCARE";
        CH1_DCOATDCFG   : string  := "DONTCARE";
        CH0_DCOBYPSATD  : string  := "DONTCARE";
        CH1_DCOBYPSATD  : string  := "DONTCARE";
        CH0_DCOSCALEI   : string  := "DONTCARE";
        CH1_DCOSCALEI   : string  := "DONTCARE";
        CH0_DCOITUNE4LSB: string  := "DONTCARE";
        CH1_DCOITUNE4LSB: string  := "DONTCARE";
        CH0_DCOIOSTUNE  : string  := "DONTCARE";
        CH1_DCOIOSTUNE  : string  := "DONTCARE";
        CH0_DCODISBDAVOID: string  := "DONTCARE";
        CH1_DCODISBDAVOID: string  := "DONTCARE";
        CH0_DCOCALDIV   : string  := "DONTCARE";
        CH1_DCOCALDIV   : string  := "DONTCARE";
        CH0_DCONUOFLSB  : string  := "DONTCARE";
        CH1_DCONUOFLSB  : string  := "DONTCARE";
        CH0_DCOIUPDNX2  : string  := "DONTCARE";
        CH1_DCOIUPDNX2  : string  := "DONTCARE";
        CH0_DCOSTEP     : string  := "DONTCARE";
        CH1_DCOSTEP     : string  := "DONTCARE";
        CH0_DCOSTARTVAL : string  := "DONTCARE";
        CH1_DCOSTARTVAL : string  := "DONTCARE";
        CH0_DCOFLTDAC   : string  := "DONTCARE";
        CH1_DCOFLTDAC   : string  := "DONTCARE";
        CH0_DCOITUNE    : string  := "DONTCARE";
        CH1_DCOITUNE    : string  := "DONTCARE";
        CH0_DCOFTNRG    : string  := "DONTCARE";
        CH1_DCOFTNRG    : string  := "DONTCARE";
        CH0_CDR_CNT4SEL : string  := "DONTCARE";
        CH1_CDR_CNT4SEL : string  := "DONTCARE";
        CH0_CDR_CNT8SEL : string  := "DONTCARE";
        CH1_CDR_CNT8SEL : string  := "DONTCARE";
        CH0_BAND_THRESHOLD: string  := "DONTCARE";
        CH1_BAND_THRESHOLD: string  := "DONTCARE";
        CH0_AUTO_FACQ_EN: string  := "DONTCARE";
        CH1_AUTO_FACQ_EN: string  := "DONTCARE";
        CH0_AUTO_CALIB_EN: string  := "DONTCARE";
        CH1_AUTO_CALIB_EN: string  := "DONTCARE";
        CH0_CALIB_CK_MODE: string  := "DONTCARE";
        CH1_CALIB_CK_MODE: string  := "DONTCARE";
        CH0_REG_BAND_OFFSET: string  := "DONTCARE";
        CH1_REG_BAND_OFFSET: string  := "DONTCARE";
        CH0_REG_BAND_SEL: string  := "DONTCARE";
        CH1_REG_BAND_SEL: string  := "DONTCARE";
        CH0_REG_IDAC_SEL: string  := "DONTCARE";
        CH1_REG_IDAC_SEL: string  := "DONTCARE";
        CH0_REG_IDAC_EN : string  := "DONTCARE";
        CH1_REG_IDAC_EN : string  := "DONTCARE";
        D_TXPLL_PWDNB   : string  := "DONTCARE";
        D_SETPLLRC      : string  := "DONTCARE";
        D_REFCK_MODE    : string  := "DONTCARE";
        D_TX_VCO_CK_DIV : string  := "DONTCARE";
        D_PLL_LOL_SET   : string  := "DONTCARE";
        D_RG_EN         : string  := "DONTCARE";
        D_RG_SET        : string  := "DONTCARE";
        D_CMUSETISCL4VCO: string  := "DONTCARE";
        D_CMUSETI4VCO   : string  := "DONTCARE";
        D_CMUSETINITVCT : string  := "DONTCARE";
        D_CMUSETZGM     : string  := "DONTCARE";
        D_CMUSETP2AGM   : string  := "DONTCARE";
        D_CMUSETP1GM    : string  := "DONTCARE";
        D_CMUSETI4CPZ   : string  := "DONTCARE";
        D_CMUSETI4CPP   : string  := "DONTCARE";
        D_CMUSETICP4Z   : string  := "DONTCARE";
        D_CMUSETICP4P   : string  := "DONTCARE";
        D_CMUSETBIASI   : string  := "DONTCARE";
        MAXLEN          : integer := 10;
        HEXLEN          : integer := 8
    );
    port(
        CH0_HDINP       : in     vl_logic;
        CH1_HDINP       : in     vl_logic;
        CH0_HDINN       : in     vl_logic;
        CH1_HDINN       : in     vl_logic;
        D_TXBIT_CLKP_FROM_ND: in     vl_logic;
        D_TXBIT_CLKN_FROM_ND: in     vl_logic;
        D_SYNC_ND       : in     vl_logic;
        D_TXPLL_LOL_FROM_ND: in     vl_logic;
        CH0_RX_REFCLK   : in     vl_logic;
        CH1_RX_REFCLK   : in     vl_logic;
        CH0_FF_RXI_CLK  : in     vl_logic;
        CH1_FF_RXI_CLK  : in     vl_logic;
        CH0_FF_TXI_CLK  : in     vl_logic;
        CH1_FF_TXI_CLK  : in     vl_logic;
        CH0_FF_EBRD_CLK : in     vl_logic;
        CH1_FF_EBRD_CLK : in     vl_logic;
        CH0_FF_TX_D_0   : in     vl_logic;
        CH1_FF_TX_D_0   : in     vl_logic;
        CH0_FF_TX_D_1   : in     vl_logic;
        CH1_FF_TX_D_1   : in     vl_logic;
        CH0_FF_TX_D_2   : in     vl_logic;
        CH1_FF_TX_D_2   : in     vl_logic;
        CH0_FF_TX_D_3   : in     vl_logic;
        CH1_FF_TX_D_3   : in     vl_logic;
        CH0_FF_TX_D_4   : in     vl_logic;
        CH1_FF_TX_D_4   : in     vl_logic;
        CH0_FF_TX_D_5   : in     vl_logic;
        CH1_FF_TX_D_5   : in     vl_logic;
        CH0_FF_TX_D_6   : in     vl_logic;
        CH1_FF_TX_D_6   : in     vl_logic;
        CH0_FF_TX_D_7   : in     vl_logic;
        CH1_FF_TX_D_7   : in     vl_logic;
        CH0_FF_TX_D_8   : in     vl_logic;
        CH1_FF_TX_D_8   : in     vl_logic;
        CH0_FF_TX_D_9   : in     vl_logic;
        CH1_FF_TX_D_9   : in     vl_logic;
        CH0_FF_TX_D_10  : in     vl_logic;
        CH1_FF_TX_D_10  : in     vl_logic;
        CH0_FF_TX_D_11  : in     vl_logic;
        CH1_FF_TX_D_11  : in     vl_logic;
        CH0_FF_TX_D_12  : in     vl_logic;
        CH1_FF_TX_D_12  : in     vl_logic;
        CH0_FF_TX_D_13  : in     vl_logic;
        CH1_FF_TX_D_13  : in     vl_logic;
        CH0_FF_TX_D_14  : in     vl_logic;
        CH1_FF_TX_D_14  : in     vl_logic;
        CH0_FF_TX_D_15  : in     vl_logic;
        CH1_FF_TX_D_15  : in     vl_logic;
        CH0_FF_TX_D_16  : in     vl_logic;
        CH1_FF_TX_D_16  : in     vl_logic;
        CH0_FF_TX_D_17  : in     vl_logic;
        CH1_FF_TX_D_17  : in     vl_logic;
        CH0_FF_TX_D_18  : in     vl_logic;
        CH1_FF_TX_D_18  : in     vl_logic;
        CH0_FF_TX_D_19  : in     vl_logic;
        CH1_FF_TX_D_19  : in     vl_logic;
        CH0_FF_TX_D_20  : in     vl_logic;
        CH1_FF_TX_D_20  : in     vl_logic;
        CH0_FF_TX_D_21  : in     vl_logic;
        CH1_FF_TX_D_21  : in     vl_logic;
        CH0_FF_TX_D_22  : in     vl_logic;
        CH1_FF_TX_D_22  : in     vl_logic;
        CH0_FF_TX_D_23  : in     vl_logic;
        CH1_FF_TX_D_23  : in     vl_logic;
        CH0_FFC_EI_EN   : in     vl_logic;
        CH1_FFC_EI_EN   : in     vl_logic;
        CH0_FFC_PCIE_DET_EN: in     vl_logic;
        CH1_FFC_PCIE_DET_EN: in     vl_logic;
        CH0_FFC_PCIE_CT : in     vl_logic;
        CH1_FFC_PCIE_CT : in     vl_logic;
        CH0_FFC_SB_INV_RX: in     vl_logic;
        CH1_FFC_SB_INV_RX: in     vl_logic;
        CH0_FFC_ENABLE_CGALIGN: in     vl_logic;
        CH1_FFC_ENABLE_CGALIGN: in     vl_logic;
        CH0_FFC_SIGNAL_DETECT: in     vl_logic;
        CH1_FFC_SIGNAL_DETECT: in     vl_logic;
        CH0_FFC_FB_LOOPBACK: in     vl_logic;
        CH1_FFC_FB_LOOPBACK: in     vl_logic;
        CH0_FFC_SB_PFIFO_LP: in     vl_logic;
        CH1_FFC_SB_PFIFO_LP: in     vl_logic;
        CH0_FFC_PFIFO_CLR: in     vl_logic;
        CH1_FFC_PFIFO_CLR: in     vl_logic;
        CH0_FFC_RATE_MODE_RX: in     vl_logic;
        CH1_FFC_RATE_MODE_RX: in     vl_logic;
        CH0_FFC_RATE_MODE_TX: in     vl_logic;
        CH1_FFC_RATE_MODE_TX: in     vl_logic;
        CH0_FFC_DIV11_MODE_RX: in     vl_logic;
        CH1_FFC_DIV11_MODE_RX: in     vl_logic;
        CH0_FFC_DIV11_MODE_TX: in     vl_logic;
        CH1_FFC_DIV11_MODE_TX: in     vl_logic;
        CH0_FFC_RX_GEAR_MODE: in     vl_logic;
        CH1_FFC_RX_GEAR_MODE: in     vl_logic;
        CH0_FFC_TX_GEAR_MODE: in     vl_logic;
        CH1_FFC_TX_GEAR_MODE: in     vl_logic;
        CH0_FFC_LDR_CORE2TX_EN: in     vl_logic;
        CH1_FFC_LDR_CORE2TX_EN: in     vl_logic;
        CH0_FFC_LANE_TX_RST: in     vl_logic;
        CH1_FFC_LANE_TX_RST: in     vl_logic;
        CH0_FFC_LANE_RX_RST: in     vl_logic;
        CH1_FFC_LANE_RX_RST: in     vl_logic;
        CH0_FFC_RRST    : in     vl_logic;
        CH1_FFC_RRST    : in     vl_logic;
        CH0_FFC_TXPWDNB : in     vl_logic;
        CH1_FFC_TXPWDNB : in     vl_logic;
        CH0_FFC_RXPWDNB : in     vl_logic;
        CH1_FFC_RXPWDNB : in     vl_logic;
        CH0_LDR_CORE2TX : in     vl_logic;
        CH1_LDR_CORE2TX : in     vl_logic;
        D_SCIWDATA0     : in     vl_logic;
        D_SCIWDATA1     : in     vl_logic;
        D_SCIWDATA2     : in     vl_logic;
        D_SCIWDATA3     : in     vl_logic;
        D_SCIWDATA4     : in     vl_logic;
        D_SCIWDATA5     : in     vl_logic;
        D_SCIWDATA6     : in     vl_logic;
        D_SCIWDATA7     : in     vl_logic;
        D_SCIADDR0      : in     vl_logic;
        D_SCIADDR1      : in     vl_logic;
        D_SCIADDR2      : in     vl_logic;
        D_SCIADDR3      : in     vl_logic;
        D_SCIADDR4      : in     vl_logic;
        D_SCIADDR5      : in     vl_logic;
        D_SCIENAUX      : in     vl_logic;
        D_SCISELAUX     : in     vl_logic;
        CH0_SCIEN       : in     vl_logic;
        CH1_SCIEN       : in     vl_logic;
        CH0_SCISEL      : in     vl_logic;
        CH1_SCISEL      : in     vl_logic;
        D_SCIRD         : in     vl_logic;
        D_SCIWSTN       : in     vl_logic;
        D_CYAWSTN       : in     vl_logic;
        D_FFC_SYNC_TOGGLE: in     vl_logic;
        D_FFC_DUAL_RST  : in     vl_logic;
        D_FFC_MACRO_RST : in     vl_logic;
        D_FFC_MACROPDB  : in     vl_logic;
        D_FFC_TRST      : in     vl_logic;
        CH0_FFC_CDR_EN_BITSLIP: in     vl_logic;
        CH1_FFC_CDR_EN_BITSLIP: in     vl_logic;
        D_SCAN_ENABLE   : in     vl_logic;
        D_SCAN_IN_0     : in     vl_logic;
        D_SCAN_IN_1     : in     vl_logic;
        D_SCAN_IN_2     : in     vl_logic;
        D_SCAN_IN_3     : in     vl_logic;
        D_SCAN_IN_4     : in     vl_logic;
        D_SCAN_IN_5     : in     vl_logic;
        D_SCAN_IN_6     : in     vl_logic;
        D_SCAN_IN_7     : in     vl_logic;
        D_SCAN_MODE     : in     vl_logic;
        D_SCAN_RESET    : in     vl_logic;
        D_CIN0          : in     vl_logic;
        D_CIN1          : in     vl_logic;
        D_CIN2          : in     vl_logic;
        D_CIN3          : in     vl_logic;
        D_CIN4          : in     vl_logic;
        D_CIN5          : in     vl_logic;
        D_CIN6          : in     vl_logic;
        D_CIN7          : in     vl_logic;
        D_CIN8          : in     vl_logic;
        D_CIN9          : in     vl_logic;
        D_CIN10         : in     vl_logic;
        D_CIN11         : in     vl_logic;
        CH0_HDOUTP      : out    vl_logic;
        CH1_HDOUTP      : out    vl_logic;
        CH0_HDOUTN      : out    vl_logic;
        CH1_HDOUTN      : out    vl_logic;
        D_TXBIT_CLKP_TO_ND: out    vl_logic;
        D_TXBIT_CLKN_TO_ND: out    vl_logic;
        D_SYNC_PULSE2ND : out    vl_logic;
        D_TXPLL_LOL_TO_ND: out    vl_logic;
        CH0_FF_RX_F_CLK : out    vl_logic;
        CH1_FF_RX_F_CLK : out    vl_logic;
        CH0_FF_RX_H_CLK : out    vl_logic;
        CH1_FF_RX_H_CLK : out    vl_logic;
        CH0_FF_TX_F_CLK : out    vl_logic;
        CH1_FF_TX_F_CLK : out    vl_logic;
        CH0_FF_TX_H_CLK : out    vl_logic;
        CH1_FF_TX_H_CLK : out    vl_logic;
        CH0_FF_RX_PCLK  : out    vl_logic;
        CH1_FF_RX_PCLK  : out    vl_logic;
        CH0_FF_TX_PCLK  : out    vl_logic;
        CH1_FF_TX_PCLK  : out    vl_logic;
        CH0_FF_RX_D_0   : out    vl_logic;
        CH1_FF_RX_D_0   : out    vl_logic;
        CH0_FF_RX_D_1   : out    vl_logic;
        CH1_FF_RX_D_1   : out    vl_logic;
        CH0_FF_RX_D_2   : out    vl_logic;
        CH1_FF_RX_D_2   : out    vl_logic;
        CH0_FF_RX_D_3   : out    vl_logic;
        CH1_FF_RX_D_3   : out    vl_logic;
        CH0_FF_RX_D_4   : out    vl_logic;
        CH1_FF_RX_D_4   : out    vl_logic;
        CH0_FF_RX_D_5   : out    vl_logic;
        CH1_FF_RX_D_5   : out    vl_logic;
        CH0_FF_RX_D_6   : out    vl_logic;
        CH1_FF_RX_D_6   : out    vl_logic;
        CH0_FF_RX_D_7   : out    vl_logic;
        CH1_FF_RX_D_7   : out    vl_logic;
        CH0_FF_RX_D_8   : out    vl_logic;
        CH1_FF_RX_D_8   : out    vl_logic;
        CH0_FF_RX_D_9   : out    vl_logic;
        CH1_FF_RX_D_9   : out    vl_logic;
        CH0_FF_RX_D_10  : out    vl_logic;
        CH1_FF_RX_D_10  : out    vl_logic;
        CH0_FF_RX_D_11  : out    vl_logic;
        CH1_FF_RX_D_11  : out    vl_logic;
        CH0_FF_RX_D_12  : out    vl_logic;
        CH1_FF_RX_D_12  : out    vl_logic;
        CH0_FF_RX_D_13  : out    vl_logic;
        CH1_FF_RX_D_13  : out    vl_logic;
        CH0_FF_RX_D_14  : out    vl_logic;
        CH1_FF_RX_D_14  : out    vl_logic;
        CH0_FF_RX_D_15  : out    vl_logic;
        CH1_FF_RX_D_15  : out    vl_logic;
        CH0_FF_RX_D_16  : out    vl_logic;
        CH1_FF_RX_D_16  : out    vl_logic;
        CH0_FF_RX_D_17  : out    vl_logic;
        CH1_FF_RX_D_17  : out    vl_logic;
        CH0_FF_RX_D_18  : out    vl_logic;
        CH1_FF_RX_D_18  : out    vl_logic;
        CH0_FF_RX_D_19  : out    vl_logic;
        CH1_FF_RX_D_19  : out    vl_logic;
        CH0_FF_RX_D_20  : out    vl_logic;
        CH1_FF_RX_D_20  : out    vl_logic;
        CH0_FF_RX_D_21  : out    vl_logic;
        CH1_FF_RX_D_21  : out    vl_logic;
        CH0_FF_RX_D_22  : out    vl_logic;
        CH1_FF_RX_D_22  : out    vl_logic;
        CH0_FF_RX_D_23  : out    vl_logic;
        CH1_FF_RX_D_23  : out    vl_logic;
        CH0_FFS_PCIE_DONE: out    vl_logic;
        CH1_FFS_PCIE_DONE: out    vl_logic;
        CH0_FFS_PCIE_CON: out    vl_logic;
        CH1_FFS_PCIE_CON: out    vl_logic;
        CH0_FFS_RLOS    : out    vl_logic;
        CH1_FFS_RLOS    : out    vl_logic;
        CH0_FFS_LS_SYNC_STATUS: out    vl_logic;
        CH1_FFS_LS_SYNC_STATUS: out    vl_logic;
        CH0_FFS_CC_UNDERRUN: out    vl_logic;
        CH1_FFS_CC_UNDERRUN: out    vl_logic;
        CH0_FFS_CC_OVERRUN: out    vl_logic;
        CH1_FFS_CC_OVERRUN: out    vl_logic;
        CH0_FFS_RXFBFIFO_ERROR: out    vl_logic;
        CH1_FFS_RXFBFIFO_ERROR: out    vl_logic;
        CH0_FFS_TXFBFIFO_ERROR: out    vl_logic;
        CH1_FFS_TXFBFIFO_ERROR: out    vl_logic;
        CH0_FFS_RLOL    : out    vl_logic;
        CH1_FFS_RLOL    : out    vl_logic;
        CH0_FFS_SKP_ADDED: out    vl_logic;
        CH1_FFS_SKP_ADDED: out    vl_logic;
        CH0_FFS_SKP_DELETED: out    vl_logic;
        CH1_FFS_SKP_DELETED: out    vl_logic;
        CH0_LDR_RX2CORE : out    vl_logic;
        CH1_LDR_RX2CORE : out    vl_logic;
        D_SCIRDATA0     : out    vl_logic;
        D_SCIRDATA1     : out    vl_logic;
        D_SCIRDATA2     : out    vl_logic;
        D_SCIRDATA3     : out    vl_logic;
        D_SCIRDATA4     : out    vl_logic;
        D_SCIRDATA5     : out    vl_logic;
        D_SCIRDATA6     : out    vl_logic;
        D_SCIRDATA7     : out    vl_logic;
        D_SCIINT        : out    vl_logic;
        D_SCAN_OUT_0    : out    vl_logic;
        D_SCAN_OUT_1    : out    vl_logic;
        D_SCAN_OUT_2    : out    vl_logic;
        D_SCAN_OUT_3    : out    vl_logic;
        D_SCAN_OUT_4    : out    vl_logic;
        D_SCAN_OUT_5    : out    vl_logic;
        D_SCAN_OUT_6    : out    vl_logic;
        D_SCAN_OUT_7    : out    vl_logic;
        D_COUT0         : out    vl_logic;
        D_COUT1         : out    vl_logic;
        D_COUT2         : out    vl_logic;
        D_COUT3         : out    vl_logic;
        D_COUT4         : out    vl_logic;
        D_COUT5         : out    vl_logic;
        D_COUT6         : out    vl_logic;
        D_COUT7         : out    vl_logic;
        D_COUT8         : out    vl_logic;
        D_COUT9         : out    vl_logic;
        D_COUT10        : out    vl_logic;
        D_COUT11        : out    vl_logic;
        D_COUT12        : out    vl_logic;
        D_COUT13        : out    vl_logic;
        D_COUT14        : out    vl_logic;
        D_COUT15        : out    vl_logic;
        D_COUT16        : out    vl_logic;
        D_COUT17        : out    vl_logic;
        D_COUT18        : out    vl_logic;
        D_COUT19        : out    vl_logic;
        D_REFCLKI       : in     vl_logic;
        D_FFS_PLOL      : out    vl_logic
    );
end DCUA;
