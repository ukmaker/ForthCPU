library verilog;
use verilog.vl_types.all;
entity ser_lslw2lwhs_0d is
    port(
        \out\           : out    vl_logic;
        vccq1           : inout  vl_logic;
        vccq2           : inout  vl_logic;
        vssq1           : inout  vl_logic;
        vssq2           : inout  vl_logic;
        enb             : in     vl_logic;
        \in\            : in     vl_logic
    );
end ser_lslw2lwhs_0d;
