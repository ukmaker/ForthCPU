library verilog;
use verilog.vl_types.all;
entity POSCDAC_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end POSCDAC_UDP;
