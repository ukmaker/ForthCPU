library verilog;
use verilog.vl_types.all;
entity NP_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end NP_UDP;
