library verilog;
use verilog.vl_types.all;
entity flash_qual is
    port(
        fl_prog_ucode_exec: out    vl_logic;
        fl_erase_exec   : out    vl_logic;
        fl_prog_done_exec: out    vl_logic;
        fl_prog_sec_exec: out    vl_logic;
        fl_prog_secplus_exec: out    vl_logic;
        fl_prog_incr_nv_exec: out    vl_logic;
        fl_prog_pwd_exec: out    vl_logic;
        fl_prog_cipher_key_exec: out    vl_logic;
        fl_prog_feature_exec: out    vl_logic;
        fl_prog_feabits_exec: out    vl_logic;
        fl_prog_otps_exec: out    vl_logic;
        fl_read_incr_nv_exec: out    vl_logic;
        fl_prog_pes_exec: out    vl_logic;
        fl_prog_mes_exec: out    vl_logic;
        fl_prog_hes_exec: out    vl_logic;
        fl_prog_trim_exec: out    vl_logic;
        fl_read_hes_exec: out    vl_logic;
        fl_init_addr_cfg_exec: out    vl_logic;
        fl_init_addr_ufm_exec: out    vl_logic;
        fl_write_addr_exec: out    vl_logic;
        fl_erase_tag_exec: out    vl_logic;
        fl_prog_tag_exec: out    vl_logic;
        fl_read_tag_exec: out    vl_logic;
        fl_mtest_exec   : out    vl_logic;
        busy_flash      : in     vl_logic;
        fea_exec_en     : in     vl_logic;
        access_sudo     : in     vl_logic;
        fl_prog_ucode_qual: in     vl_logic;
        fl_erase_qual   : in     vl_logic;
        fl_prog_done_qual: in     vl_logic;
        fl_prog_sec_qual: in     vl_logic;
        fl_prog_secplus_qual: in     vl_logic;
        fl_init_addr_qual: in     vl_logic;
        fl_write_addr_qual: in     vl_logic;
        fl_prog_incr_nv_qual: in     vl_logic;
        fl_read_incr_nv_qual: in     vl_logic;
        fl_prog_password_qual: in     vl_logic;
        fl_prog_cipher_key_qual: in     vl_logic;
        fl_prog_feature_qual: in     vl_logic;
        fl_prog_feabits_qual: in     vl_logic;
        fl_prog_otps_qual: in     vl_logic;
        fl_init_addr_ufm_qual: in     vl_logic;
        fl_prog_tag_qual: in     vl_logic;
        fl_erase_tag_qual: in     vl_logic;
        fl_read_tag_qual: in     vl_logic;
        fl_prog_pes_qual: in     vl_logic;
        fl_prog_mes_qual: in     vl_logic;
        fl_prog_hes_qual: in     vl_logic;
        fl_prog_trim_qual: in     vl_logic;
        fl_read_hes_qual: in     vl_logic;
        fl_mtest_qual   : in     vl_logic
    );
end flash_qual;
