library verilog;
use verilog.vl_types.all;
entity hsc_sbnx16v1e is
    port(
        A               : in     vl_logic;
        Z               : out    vl_logic
    );
end hsc_sbnx16v1e;
