library verilog;
use verilog.vl_types.all;
entity TGM2_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end TGM2_UDP;
