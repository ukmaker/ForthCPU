library verilog;
use verilog.vl_types.all;
entity config_io is
    port(
        pi_scl_d        : out    vl_logic;
        pi_sda_d        : out    vl_logic;
        shbsrn          : out    vl_logic;
        pll_mfg_ts      : out    vl_logic_vector(1 downto 0);
        pll_mfg_md_n    : out    vl_logic_vector(1 downto 0);
        bsmode          : out    vl_logic;
        intest          : out    vl_logic;
        ts_all          : out    vl_logic;
        cib_i2c_sclen   : out    vl_logic;
        cib_i2c_sdaen   : out    vl_logic;
        jtagenb_pin     : out    vl_logic;
        done_pin        : out    vl_logic;
        initn_pin       : out    vl_logic;
        programn_pin    : out    vl_logic;
        tck_pin         : out    vl_logic;
        tms_pin         : out    vl_logic;
        cib_mspi_csn    : out    vl_logic_vector(7 downto 1);
        csspin          : out    vl_logic;
        program_md_n    : out    vl_logic;
        done_md_n       : out    vl_logic;
        done_ts         : out    vl_logic;
        init_md_n       : out    vl_logic;
        init_ts         : out    vl_logic;
        mspi_md_n       : out    vl_logic;
        mclk_out        : out    vl_logic;
        mclk_ts         : out    vl_logic;
        i2c_md_n        : out    vl_logic;
        scl             : out    vl_logic;
        sda             : out    vl_logic;
        scl_ts          : out    vl_logic;
        sda_ts          : out    vl_logic;
        si              : out    vl_logic;
        si_md_n         : out    vl_logic;
        si_ts           : out    vl_logic;
        so              : out    vl_logic;
        so_md_n         : out    vl_logic;
        so_ts           : out    vl_logic;
        jtag_md_n       : out    vl_logic;
        tdo_ts          : out    vl_logic;
        pi_scl          : in     vl_logic;
        pi_sda          : in     vl_logic;
        mfg_pll_out     : in     vl_logic_vector(1 downto 0);
        shiftdr_bs      : in     vl_logic;
        progn_persist   : in     vl_logic;
        initn_persist   : in     vl_logic;
        donep_persist   : in     vl_logic;
        cib_i2c_scle    : in     vl_logic;
        cib_i2c_sdae    : in     vl_logic;
        mc1_mspi_persist: in     vl_logic;
        mc1_sspi_persist: in     vl_logic;
        mclk_o_2nd      : in     vl_logic;
        mclk_oe_2nd     : in     vl_logic;
        miso_o_2nd      : in     vl_logic;
        miso_oe_2nd     : in     vl_logic;
        mosi_o_2nd      : in     vl_logic;
        mosi_oe_2nd     : in     vl_logic;
        jtagenb         : in     vl_logic;
        donein          : in     vl_logic;
        initin_n        : in     vl_logic;
        programn        : in     vl_logic;
        bsmode1         : in     vl_logic;
        bsmode2         : in     vl_logic;
        bsmode3         : in     vl_logic;
        tck             : in     vl_logic;
        tms             : in     vl_logic;
        mcsn_o          : in     vl_logic_vector(7 downto 0);
        mcsn_oe         : in     vl_logic_vector(7 downto 0);
        mcsn_o_cib      : in     vl_logic_vector(7 downto 0);
        mcsn_oe_cib     : in     vl_logic_vector(7 downto 0);
        done_goe        : in     vl_logic;
        data_o          : in     vl_logic_vector(3 downto 0);
        data_oe         : in     vl_logic_vector(3 downto 0);
        mclk_o          : in     vl_logic;
        mclk_oe         : in     vl_logic;
        jtag_persist    : in     vl_logic;
        tdo_oe          : in     vl_logic;
        donep_oe        : in     vl_logic;
        initn_oe        : in     vl_logic;
        sspi_oe         : in     vl_logic;
        sspi_so         : in     vl_logic;
        sda_oe_pad      : in     vl_logic;
        scl_oe_pad      : in     vl_logic;
        sda_out_pad     : in     vl_logic;
        scl_out_pad     : in     vl_logic
    );
end config_io;
