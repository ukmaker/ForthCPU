library verilog;
use verilog.vl_types.all;
entity pcs_inv_6 is
    port(
        A               : in     vl_logic;
        X               : out    vl_logic
    );
end pcs_inv_6;
