library verilog;
use verilog.vl_types.all;
entity pcs_ch_dp is
    port(
        bus8bit_sel     : in     vl_logic;
        txp_clk         : in     vl_logic;
        rstb_txp        : in     vl_logic;
        rxr_clk         : in     vl_logic;
        rstb_rxr        : in     vl_logic;
        ebrd_clk        : in     vl_logic;
        rstb_ebrd       : in     vl_logic;
        fbw_clk         : in     vl_logic;
        rstb_fbw        : in     vl_logic;
        txf_clk         : in     vl_logic;
        rstb_txf        : in     vl_logic;
        rxf_clk         : in     vl_logic;
        rstb_rxf        : in     vl_logic;
        txd_fifo_lb     : in     vl_logic_vector(9 downto 0);
        serdes_rxd      : in     vl_logic_vector(9 downto 0);
        txd_sd          : out    vl_logic_vector(9 downto 0);
        tobist_data     : out    vl_logic_vector(9 downto 0);
        bist_rx_data_sel: in     vl_logic;
        fmbist_data     : in     vl_logic_vector(9 downto 0);
        ff_tx_d         : in     vl_logic_vector(23 downto 0);
        ff_rx_d         : out    vl_logic_vector(23 downto 0);
        plol            : in     vl_logic;
        pcie_txdetrx_pr2tlb: in     vl_logic;
        pcie_txcomp     : in     vl_logic;
        pcie_txeleci    : in     vl_logic;
        pcie_rxpolarity : in     vl_logic;
        pcie_powerdown  : in     vl_logic_vector(1 downto 0);
        pcie_p2         : out    vl_logic;
        phystatus       : out    vl_logic;
        ffc_pcie_ct     : in     vl_logic;
        pcie_cts        : out    vl_logic;
        ffc_pcie_det_en : in     vl_logic;
        pci_det_en      : out    vl_logic;
        ffc_signal_detect: in     vl_logic;
        ffc_enable_cgalign: in     vl_logic;
        ffc_fb_loopback : in     vl_logic;
        ffc_sb_pfifo_lp : in     vl_logic;
        ffc_sb_inv_rx   : in     vl_logic;
        ffc_cdr_en_bitslip: in     vl_logic;
        ffs_ls_sync_status: out    vl_logic;
        ffs_cc_overrun  : out    vl_logic;
        ffs_cc_underrun : out    vl_logic;
        ffs_rxfbfifo_error: out    vl_logic;
        ffs_txfbfifo_error: out    vl_logic;
        pcie_det_done   : in     vl_logic;
        pci_connect     : in     vl_logic;
        ffc_ei_en       : in     vl_logic;
        pci_ei_en       : out    vl_logic;
        pcie_det_time_sel: out    vl_logic_vector(1 downto 0);
        rx_ch           : out    vl_logic;
        char_test_data  : in     vl_logic_vector(9 downto 0);
        char_test_mode  : in     vl_logic;
        pfifo_error     : in     vl_logic;
        prbs_error      : out    vl_logic;
        pcs_ctl_2_ch_01 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_3_ch_02 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_4_ch_03 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_5_ch_04 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_6_ch_05 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_7_ch_06 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_8_ch_07 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_9_ch_08 : in     vl_logic_vector(7 downto 0);
        pcs_ctl_10_ch_09: in     vl_logic_vector(7 downto 0);
        pcs_ctl_11_ch_0a: in     vl_logic_vector(7 downto 0);
        pcs_ctl_12_ch_0b: in     vl_logic_vector(7 downto 0);
        pcs_ctl_13_ch_0c: in     vl_logic_vector(7 downto 0);
        pcs_ctl_14_ch_0d: in     vl_logic_vector(7 downto 0);
        pcs_ctl_15_ch_0e: in     vl_logic_vector(7 downto 0);
        pcs_sts_1_ch_20 : out    vl_logic_vector(7 downto 0);
        pcs_sts_3_ch_22 : out    vl_logic_vector(7 downto 0);
        pcs_sts_5_ch_24 : out    vl_logic_vector(7 downto 0);
        pcs_sts_6_ch_25 : out    vl_logic_vector(7 downto 0);
        uc_mode         : in     vl_logic;
        fc_mode         : in     vl_logic;
        pcie_mode       : in     vl_logic;
        rio_mode        : in     vl_logic;
        wa_mode         : in     vl_logic;
        xge_mode        : in     vl_logic;
        lsm_eca         : in     vl_logic;
        pcs_ctl_3_dl_02 : in     vl_logic_vector(7 downto 0);
        cdr_en_bitslip  : out    vl_logic
    );
end pcs_ch_dp;
