library verilog;
use verilog.vl_types.all;
entity faultlog_prgm is
    generic(
        st_reset        : integer := 0;
        st_findrow1     : integer := 1;
        st_findrow2     : integer := 3;
        st_findrow3     : integer := 2;
        st_findrow4     : integer := 6;
        st_findrow5     : integer := 7;
        st_findrow6     : integer := 5;
        st_detect0      : integer := 4;
        st_detect1      : integer := 12;
        st_setupa       : integer := 13;
        st_setup        : integer := 15;
        st_soft1        : integer := 14;
        st_soft2        : integer := 10;
        st_hard1        : integer := 11;
        st_cancel1      : integer := 9;
        st_cancel2      : integer := 8;
        st_prgm_setup1  : integer := 24;
        st_prgm_setup2  : integer := 16;
        st_prgm_eep     : integer := 17;
        st_finish1      : integer := 19;
        st_finish2      : integer := 18;
        st_finish3      : integer := 22
    );
    port(
        mc_twifl_data   : out    vl_logic_vector(7 downto 0);
        faultlog_sel_3wi: out    vl_logic;
        flut_col_addr   : out    vl_logic_vector(2 downto 0);
        flut_row_addr   : out    vl_logic_vector(3 downto 0);
        flut_load_datareg: out    vl_logic;
        faultlog_load_soft_datareg: out    vl_logic;
        force_erasprgm_st3: out    vl_logic;
        twi_fl_prgm_eep : out    vl_logic;
        faultlog_in_progress: out    vl_logic;
        clear_verrdall_iflg: out    vl_logic;
        clear_rdsoftfault_iflg: out    vl_logic;
        faultlog_full   : out    vl_logic;
        eep_shdw_ready  : out    vl_logic;
        examine_fldonebit: out    vl_logic;
        faultlog_next_row: out    vl_logic_vector(3 downto 0);
        flrden_stat     : out    vl_logic_vector(7 downto 0);
        flclr_ep_iflgs  : out    vl_logic;
        rst_erase_prgm_stmach: out    vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        refresh_on      : in     vl_logic;
        usertag_enable  : in     vl_logic;
        mc_mcb_in       : in     vl_logic_vector(7 downto 0);
        twi_start       : in     vl_logic;
        twi_rdat_read   : in     vl_logic;
        twi_rdat_data_from_latch: in     vl_logic_vector(7 downto 0);
        twi_flid_shdw   : in     vl_logic_vector(7 downto 0);
        twi_fl_record   : in     vl_logic;
        twi_fl_soft     : in     vl_logic;
        ld_wr_data_reg  : in     vl_logic;
        writeusertag_iflg: in     vl_logic;
        flut_reset_flutaddrregctr: in     vl_logic;
        flut_incr_flutaddrregupctr: in     vl_logic;
        erase_prgrm_active: in     vl_logic;
        eraseflut_iflg  : in     vl_logic;
        flut_load_flutaddrregupctr: in     vl_logic;
        not_verrdall_iflg: in     vl_logic;
        not_rdsoftfault : in     vl_logic;
        rdusertag_iflg  : in     vl_logic;
        incr_rd_addr_ctr: in     vl_logic;
        verfault_iflg   : in     vl_logic;
        load_rdfaultenlat: in     vl_logic;
        fault_i2csa_erasprgm_iflg: in     vl_logic
    );
end faultlog_prgm;
