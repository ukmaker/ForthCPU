library verilog;
use verilog.vl_types.all;
entity LN4_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end LN4_UDP;
