library verilog;
use verilog.vl_types.all;
entity njtag_cmd_dec is
    port(
        bypass_c        : out    vl_logic;
        verify_id_c     : out    vl_logic;
        idcode_pub_c    : out    vl_logic;
        uidcode_pub_c   : out    vl_logic;
        usercode_c      : out    vl_logic;
        read_temp_c     : out    vl_logic;
        lsc_device_ctrl_c: out    vl_logic;
        lsc_shift_password_c: out    vl_logic;
        lsc_read_status_c: out    vl_logic;
        lsc_check_busy_c: out    vl_logic;
        lsc_refresh_c   : out    vl_logic;
        lsc_bitstream_burst_c: out    vl_logic;
        lsc_i2ci_crbr_wt_c: out    vl_logic;
        lsc_i2ci_txdr_wt_c: out    vl_logic;
        lsc_i2ci_rxdr_rd_c: out    vl_logic;
        lsc_i2ci_sr_rd_c: out    vl_logic;
        lsc_prog_spi_c  : out    vl_logic;
        idcode_prv_c    : out    vl_logic;
        read_pes_c      : out    vl_logic;
        isc_enable_c    : out    vl_logic;
        isc_enable_x_c  : out    vl_logic;
        isc_disable_c   : out    vl_logic;
        isc_program_c   : out    vl_logic;
        isc_noop_c      : out    vl_logic;
        isc_prog_ucode_c: out    vl_logic;
        isc_read_c      : out    vl_logic;
        isc_erase_c     : out    vl_logic;
        isc_prog_done_c : out    vl_logic;
        isc_erase_done_c: out    vl_logic;
        isc_prog_sec_c  : out    vl_logic;
        isc_prog_secplus_c: out    vl_logic;
        isc_data_shift_c: out    vl_logic;
        isc_addr_shift_c: out    vl_logic;
        lsc_init_addr_c : out    vl_logic;
        lsc_write_addr_c: out    vl_logic;
        lsc_prog_incr_rti_c: out    vl_logic;
        lsc_prog_incr_enc_c: out    vl_logic;
        lsc_prog_incr_cmp_c: out    vl_logic;
        lsc_prog_incr_cne_c: out    vl_logic;
        lsc_vfy_incr_rti_c: out    vl_logic;
        lsc_prog_ctrl0_c: out    vl_logic;
        lsc_read_ctrl0_c: out    vl_logic;
        lsc_reset_crc_c : out    vl_logic;
        lsc_read_crc_c  : out    vl_logic;
        lsc_prog_sed_crc_c: out    vl_logic;
        lsc_read_sed_crc_c: out    vl_logic;
        lsc_prog_password_c: out    vl_logic;
        lsc_read_password_c: out    vl_logic;
        lsc_prog_cipher_key_c: out    vl_logic;
        lsc_read_cipher_key_c: out    vl_logic;
        lsc_prog_feature_c: out    vl_logic;
        lsc_read_feature_c: out    vl_logic;
        lsc_prog_feabits_c: out    vl_logic;
        lsc_read_feabits_c: out    vl_logic;
        lsc_prog_otps_c : out    vl_logic;
        lsc_read_otps_c : out    vl_logic;
        lsc_write_comp_dic_c: out    vl_logic;
        lsc_write_bus_addr_c: out    vl_logic;
        lsc_pcs_write_c : out    vl_logic;
        lsc_pcs_read_c  : out    vl_logic;
        lsc_ebr_write_c : out    vl_logic;
        lsc_ebr_read_c  : out    vl_logic;
        lsc_prog_incr_nv_c: out    vl_logic;
        lsc_read_incr_nv_c: out    vl_logic;
        lsc_init_addr_ufm_c: out    vl_logic;
        lsc_prog_tag_c  : out    vl_logic;
        lsc_erase_tag_c : out    vl_logic;
        lsc_read_tag_c  : out    vl_logic;
        lsc_chip_select_c: out    vl_logic;
        lsc_flow_through_c: out    vl_logic;
        lsc_jump_c      : out    vl_logic;
        nj_invalid_c    : out    vl_logic;
        njcommand       : in     vl_logic_vector(7 downto 0)
    );
end njtag_cmd_dec;
