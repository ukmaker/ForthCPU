library verilog;
use verilog.vl_types.all;
entity ser_tx_misc is
    port(
        bit_from_nd_eno : out    vl_logic;
        bs2pado         : out    vl_logic;
        irefpwdnbo      : out    vl_logic;
        ldr_core2tx_selo: out    vl_logic;
        ldr_core2txo    : out    vl_logic;
        pci_connect     : out    vl_logic;
        pci_connect_sts : out    vl_logic;
        pci_det_cto     : out    vl_logic;
        pci_det_done    : out    vl_logic;
        pci_det_eno     : out    vl_logic;
        pci_ei_eno      : out    vl_logic;
        pcie_modeo      : out    vl_logic;
        rate_mode_txo   : out    vl_logic;
        rterm_txo       : out    vl_logic_vector(3 downto 0);
        sync_local_eno  : out    vl_logic;
        sync_nd_eno     : out    vl_logic;
        tck             : out    vl_logic;
        tdo             : out    vl_logic_vector(9 downto 0);
        tdrv_dat_selo   : out    vl_logic_vector(1 downto 0);
        tdrv_post_eno   : out    vl_logic;
        tdrv_pre_eno    : out    vl_logic;
        tdrv_slice0_curo: out    vl_logic_vector(2 downto 0);
        tdrv_slice0_selo: out    vl_logic_vector(1 downto 0);
        tdrv_slice1_curo: out    vl_logic_vector(2 downto 0);
        tdrv_slice1_selo: out    vl_logic_vector(1 downto 0);
        tdrv_slice2_curo: out    vl_logic_vector(1 downto 0);
        tdrv_slice2_selo: out    vl_logic_vector(1 downto 0);
        tdrv_slice3_curo: out    vl_logic_vector(1 downto 0);
        tdrv_slice3_selo: out    vl_logic_vector(1 downto 0);
        tdrv_slice4_curo: out    vl_logic;
        tdrv_slice4_selo: out    vl_logic_vector(1 downto 0);
        tdrv_slice5_curo: out    vl_logic;
        tdrv_slice5_selo: out    vl_logic_vector(1 downto 0);
        tpwdnbo         : out    vl_logic;
        tx_bs_modeo     : out    vl_logic;
        tx_cm_selo      : out    vl_logic_vector(1 downto 0);
        tx_div11_selo   : out    vl_logic;
        tx_post_signo   : out    vl_logic;
        tx_pre_signo    : out    vl_logic;
        vcc             : inout  vl_logic;
        vccatx          : inout  vl_logic;
        vss             : inout  vl_logic;
        vssatx          : inout  vl_logic;
        vssatxs         : inout  vl_logic;
        bit_from_nd_en  : in     vl_logic;
        bs2pad          : in     vl_logic;
        ldr_core2tx     : in     vl_logic;
        ldr_core2tx_sel : in     vl_logic;
        macropdb        : in     vl_logic;
        pci_connectin   : in     vl_logic;
        pci_det_ct      : in     vl_logic;
        pci_det_donein  : in     vl_logic;
        pci_det_en      : in     vl_logic;
        pci_ei_en       : in     vl_logic;
        pcie_mode       : in     vl_logic;
        rate_mode_tx    : in     vl_logic;
        rpwdnbin        : in     vl_logic;
        rterm_tx        : in     vl_logic_vector(3 downto 0);
        rx_bs_modein    : in     vl_logic;
        sync_local_en   : in     vl_logic;
        sync_nd_en      : in     vl_logic;
        tckin           : in     vl_logic;
        td              : in     vl_logic_vector(9 downto 0);
        tdrv_dat_sel    : in     vl_logic_vector(1 downto 0);
        tdrv_post_en    : in     vl_logic;
        tdrv_pre_en     : in     vl_logic;
        tdrv_slice0_cur : in     vl_logic_vector(2 downto 0);
        tdrv_slice0_sel : in     vl_logic_vector(1 downto 0);
        tdrv_slice1_cur : in     vl_logic_vector(2 downto 0);
        tdrv_slice1_sel : in     vl_logic_vector(1 downto 0);
        tdrv_slice2_cur : in     vl_logic_vector(1 downto 0);
        tdrv_slice2_sel : in     vl_logic_vector(1 downto 0);
        tdrv_slice3_cur : in     vl_logic_vector(1 downto 0);
        tdrv_slice3_sel : in     vl_logic_vector(1 downto 0);
        tdrv_slice4_cur : in     vl_logic;
        tdrv_slice4_sel : in     vl_logic_vector(1 downto 0);
        tdrv_slice5_cur : in     vl_logic;
        tdrv_slice5_sel : in     vl_logic_vector(1 downto 0);
        tpwdnb          : in     vl_logic;
        tx_bs_mode      : in     vl_logic;
        tx_cm_sel       : in     vl_logic_vector(1 downto 0);
        tx_div11_sel    : in     vl_logic;
        tx_post_sign    : in     vl_logic;
        tx_pre_sign     : in     vl_logic
    );
end ser_tx_misc;
