library verilog;
use verilog.vl_types.all;
entity pcs_clk_rst is
    port(
        asyn_mode       : in     vl_logic;
        ff_rxi_clk      : in     vl_logic_vector(1 downto 0);
        ff_txi_clk      : in     vl_logic_vector(1 downto 0);
        ff_ebrd_clk     : in     vl_logic_vector(1 downto 0);
        rxr_clk_sd      : in     vl_logic_vector(1 downto 0);
        txp_clk_sd      : in     vl_logic_vector(1 downto 0);
        refc2core       : in     vl_logic;
        ffc_ck_core_rx  : in     vl_logic_vector(1 downto 0);
        ffc_ck_core_tx  : in     vl_logic;
        tck_aux_full    : in     vl_logic;
        cfg_clk         : in     vl_logic;
        cin             : in     vl_logic_vector(11 downto 0);
        sel_sd_rx_clk   : in     vl_logic_vector(1 downto 0);
        sel_test_clk    : in     vl_logic;
        ffc_rx_lane_rst : in     vl_logic_vector(1 downto 0);
        ffc_tx_lane_rst : in     vl_logic_vector(1 downto 0);
        ffc_dual_rst    : in     vl_logic;
        lane_rx_rst     : in     vl_logic_vector(1 downto 0);
        lane_tx_rst     : in     vl_logic_vector(1 downto 0);
        ff_tx_f_clk_dis : in     vl_logic_vector(1 downto 0);
        ff_tx_h_clk_en  : in     vl_logic_vector(1 downto 0);
        ff_rx_f_clk_dis : in     vl_logic_vector(1 downto 0);
        ff_rx_h_clk_en  : in     vl_logic_vector(1 downto 0);
        bist_rpt_ch_sel : in     vl_logic;
        bist_en         : in     vl_logic;
        char_mode       : in     vl_logic;
        rst_ctl_1_dl_10 : in     vl_logic_vector(2 downto 0);
        ffc_macro_rst   : in     vl_logic;
        ffc_trst        : in     vl_logic;
        ffc_rrst        : in     vl_logic_vector(1 downto 0);
        rrst_reg        : in     vl_logic_vector(1 downto 0);
        ffc_pfifo_clr   : in     vl_logic_vector(1 downto 0);
        full_d          : in     vl_logic_vector(1 downto 0);
        empty_d         : in     vl_logic_vector(1 downto 0);
        plol            : in     vl_logic;
        txpll_lol_from_nd: in     vl_logic;
        pcs_ctl_3_ch_02_710: in     vl_logic_vector(3 downto 0);
        pcs_ctl_3_ch_02_32: in     vl_logic_vector(3 downto 0);
        sciwstn         : in     vl_logic;
        scan_enable     : in     vl_logic;
        scan_in_7       : in     vl_logic;
        done_cfg        : in     vl_logic;
        disable_dcu     : in     vl_logic;
        txp_clk         : out    vl_logic_vector(1 downto 0);
        txf_clk         : out    vl_logic_vector(1 downto 0);
        rxr_clk         : out    vl_logic_vector(1 downto 0);
        ebrd_clk        : out    vl_logic_vector(1 downto 0);
        fbw_clk         : out    vl_logic_vector(1 downto 0);
        rxf_clk         : out    vl_logic_vector(1 downto 0);
        ff_rx_f_clk     : out    vl_logic_vector(1 downto 0);
        ff_rx_h_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_f_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_h_clk     : out    vl_logic_vector(1 downto 0);
        ff_tx_pclk      : out    vl_logic_vector(1 downto 0);
        ff_rx_pclk      : out    vl_logic_vector(1 downto 0);
        refck2core      : out    vl_logic;
        ck_core_rx      : out    vl_logic_vector(1 downto 0);
        ck_core_tx      : out    vl_logic;
        bist_tx_clk     : out    vl_logic;
        bist_rx_clk     : out    vl_logic;
        bist_wrst       : out    vl_logic;
        bist_rrst       : out    vl_logic;
        reg_load        : out    vl_logic;
        goe_r2          : out    vl_logic;
        goe_load        : out    vl_logic;
        cout_19         : out    vl_logic;
        cout_16         : out    vl_logic;
        cout_2          : out    vl_logic;
        cout_0          : out    vl_logic;
        rstb_txf        : out    vl_logic_vector(1 downto 0);
        rstb_txp        : out    vl_logic_vector(1 downto 0);
        rstb_ebrd       : out    vl_logic_vector(1 downto 0);
        rstb_rxr        : out    vl_logic_vector(1 downto 0);
        rstb_fbw        : out    vl_logic_vector(1 downto 0);
        rstb_rxf        : out    vl_logic_vector(1 downto 0);
        macrorst        : out    vl_logic;
        trst            : out    vl_logic;
        rrst            : out    vl_logic_vector(1 downto 0);
        pfifow_clr      : out    vl_logic_vector(1 downto 0);
        pfifor_clr      : out    vl_logic_vector(1 downto 0);
        txpll_lol_to_nd : out    vl_logic;
        char_test_data  : out    vl_logic_vector(9 downto 0);
        char_test_mode  : out    vl_logic;
        cib_dis         : out    vl_logic
    );
end pcs_clk_rst;
