`include "../../constants.v"

/*****************************************
* 
*****************************************/
module instructionLatch(
	
	
);



endmodule